// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GlqWlhot5+LrPLGJF2NIWN0CR3PxXj4VNjbYjbJtDJzavNPoUUCpDnURhVq/6XUK
/aBKoo8gaVvXrDT1B/O/huLupDtv0xcJjzOOT3z3aKMVj94fBRbZ5YsEGqhTnycb
lRKR+fRgBUy3U8NHK+Ho0kbVhw2oeOxxX8xIVrhLa5g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11456)
lxS/ucoS9AuTKkuiZQABrhPu2DL7EvynLmVvwdZyZG/XHMz4hSuAlwPDw9sZ4YIe
zOsNvUhmZrvefYyH4Fu9xQzi8fyNOqJ1Y97I2PQ3VSTotzmOvgXKin+B6G98gTQV
zUvTNIR5qGN0vTuO5WA+ixD+mxh/qDay6t/wHvOanFU6bQFe9+FQoGM8D3/U5h1g
81ZKRgZSYLZvBDELh3GokHu3YX1YwM+6mYTUSpCtV7hOi8tJBMmWTCLv334nRsEz
1XapX4Mthzs/QQyovFlHJUvAARcyC1PQHGZKVerpvQJlElfXJwqlLxVDBGeJVcLW
sxu9w/2v0PCd9tDxRpFrr7uHTFuXf+KwwUwN1V+OC3/00k0Uxi8/EKPBJPxSbuNV
hEe9I/IRnBNq6LY/A0d3ke/NHAVovfoSFMAOdWW1TzSR+0ZobirxkfFBauYOGDpd
nDFY6pCrHDxdKWknjbznkAPMv0e/iNfrGGhxIUO6XRNluiUwXIfK3bqRughGn7ZD
KMhD6qmU+QFQvkkrEeqJx1IB7gAFpgTRHJkMEI8+sLufHK5WO+gSnKq0Ad2NlgTy
8UhEM3zEmFEO5nXoyNTMzfBvlF/jRzMBmMkij2bFe08Nx74rkU4dpwxG34KlYYv5
3e8/e4K7kVVeECcG0VFj29+WBllosZg3pFTMrXnM15snwGP1qOAMCeyNxLsNOrtZ
UhwVd8lsNXvWSpDogGF7vA7fwoElbuEqrD/c83dgy1UozUBGrhnBcM3JjL87z3uj
R4z7BLkP7NqiMt2GB0EEHUzD9IFfAv4HOGcUMoCnIQitrgv43UIciUnKcNBKSM/1
7MznL5xIoP+TSlVam5n5vHVpRkXTJeXh4Yb5Pk3XfrFutsSVyL90KuobLNlrLvJA
wDJgms2PDHj5KvOBcGXoeOkCzB05/2dQ68lyKq/fS+zsK33S2uTki6x/3wRjT/fd
MbZVDw/R11iLFRwjRzmBrSFEkepD+f3XUg8M7h7qJbgYdX+K8JNjQbU/lfitmtpZ
8gJvNPTpwSq12a5cVn3QCqh5jFRiiv1CXdnV3Np52sAxxufAzZne5luqMr+I0cYa
q9K89Po8f54Q8b8/vbCPJ8JyRC6/nRRw3nBELTqHgRRGQh+Mxld3pCFiyItK+T99
S7QiYQK/EifkkwVWynFbLxOsNyGqr5oGcaQHq1jOxFbBCQtTGb3alclMQlegf3PB
S0jdmLbFMOR2A8PmlBJ6HoNHZLS89mAOPvrZYqEFR2ccLqSu62WPgIdiuhYDxPry
JrJ5wvjPO2gUvWbgG7RMlFNHnUmsbau+PKbDH9Jh8r/CAAo7uz74dFrQYk+iCjY7
7u5BuvO7YZsFnCINmKgtoA3RpKa9yy8njdP705IoCwcqUTTMNk2UaWyaPi01omGt
OuZBiZIegrONm4hU5uc1gSHiroGje9SriTfF50b9szg/4lZuP2msjzZuLVic/YIJ
X35iwyXQefkG8vtNRYWFByOrdbN5OB0kj8gB08ghrrNhGz9ayeCXYEr2tmQ9Lkxp
OwYZlV+FEfiLnlcF0p3ZFGZ5YzX7p15dYHGIqLUhvH5hVlxxE/WPVA76e8eQ/aB4
mo/RJ8byYN2mJwHYDBlSt20ZPvIdKxC0xC19po4qnIfeZvaMnotSt3HhuScEeNmh
9cw8z9i1LYQPfSpMi6SgqsLdb++ZQPdJ1nYPUFwhDXY8fDHXzLKCg1Lmts14/SHl
jbSxeRAd2e/ys9Q5fXRxcs/ABuSYH+eBf/bqxVo2NeqE/4DKftCIZJVSZDe80SZG
3czHIgtUT1i7KNDwaWpnurylhTjeDMXcOHbzQmJd6hrbVqiuqkGzYLs0ITs60uaM
+GV4KX6ZqSdiNkkl07rQB4JfaNpRR+ErDuIj0XUKp8TNIZcV1JNq1zBd+UM7Qx8x
yBENP8vFrmkyRnYSGH1zIvfsXuvFW16O4MZjKGVHUxwkCpK1CBs6RCd0jX53HQ1o
YWBvH/qKy7fXyCGqN+h3yve2gydIEwydRS+qDHcE+HWxKjauScEYLsSya+xFZZ8F
RtPEBTaIptcvC5Wlk8tlyExkan5LiquNj0E8gEiuUYW8cDKqRIP7p1WHODWpaA+q
Mo+vIMkO/dmiu0IbRTTt7KOb3jt5w9duLjPF72YWaME1kmXn7hMzgKXBXWKYDdNr
ndj05WeErANiWaERnJPTsq459VlvJRpkMYaFqUeGhkxvT9iBgSw+pdNA2u3PbzBc
DH8KgOpP6VBI0uqlQipJ0Zp6p+wFK6R59nGWTDYZLoUyDs1nUdjjWPiAVCFAMF9j
30mZ2HVZgX4mA7iM/Cj3GGmB1PF/D37VYWbnCWp/+ucTX+q34aU1j9e9R3x86sSN
FAeo9Ur+nf/faUxjVzo6KXyl3jQ2hOTWGeyGZLEfSTgbV3Id30GhFKUz94Q+vSm5
Nn7BjL2RCPWjjbwLrt+N2dPgO9cfItfo3J+Ectda9R6XOcYQgQzunaQ9N6wBg2W2
gMazrZ168+DZbf2bPqCEYqb9013nKS6jqgpuuN1w41JjJR1xZ+T35g3Fh5LxrliZ
OYYdpyOEwhnroGCEV3UeoUo4nh3PVuSGlhpf0fUg8G2/sUIYgnIP5WC9OJIPtJm1
qpznYB7WKiNWjHKZDRqzdjvOXp8l66k8lg3PX39BmCvHW1VrTOFoIEzPr/PAoSVO
OJvnZ09G+jppiX0ST78rksdyvQ7KghC6L1zv2Hpl/vZWa1el1pEGa7vA5y7s7aVN
rBAFZoCc1M97iDCuRbfJpGenRqFdUXAvKAX5PKBPyi1sMOpy3BYEcwCzjd6f5XDk
uIVT4g8SdS2nFlf4HFGx4fmGdtliwgPURc5Gk8eKDtfRL9BeoZy9aNSr6C4dIZNe
Bi8KdaQWO4E5gjCpJRVGKZebzsZKsEC5xfEyZCN+5wBp3Dpdbl9N3s20x6oTxe7A
Tsv5fmtU2RLpJXdhp0n5vHiF75B+FwAtBoLhEEDgN19lskvktFV4f7iOI0yvO0Pg
sGvCoJh1x1TD0tH655/zsCFYLj66H0jnwGHWacKExy0YwLF0dKSrFbt1bTZY3n+b
spPPJmufpyrIpw/4DpmQ1izm7Y9p5KevZBkyUUHKlpTUQv4Wa9pPHuHcvbc/nMaL
BG7zJr6y/gCLFgKijJZi87L7AsgBUuoqMTGd5HIqz3VxTpfjcK82mxTVSCdHpUNi
OysUuEcefusTcWre54YlQNHO+y1zWy5RMusqiTMY6SJrK9+HMsLWDOOjZX8cbycg
C39SN14KaKvpICUwZFqJEPC/E2DTUkia80dztG/7Qfr/F8YqrsXyKxDbv1uUTP7K
u+I5umh5diF6U7VwAgDpIYwuRba66OtNxyIjZDPUd/Fj5y9YoF9U5iQzYqjTGqOw
Lb6n1HgtovqAqNkevSMXoTNHxFgLkmWWq3PkGibHgCEjAhmyhrDxumRA9bSQlXG5
N7XwL0X8syacTFy7JP20PLGbjS/2x++EerRCUH2ffyU9ZexdHSMZfzec9DmWMSac
LC9eoLb9Q+rZ7mzDtFaDHBTlcqwmGxLsDvJoH5i7lg4YUSJQ5NzBRAFxNjx1UlPQ
tDn7V1iek8M/G+xuXZDpEPYvLy4KowHy3gMeu4pyGsg2wX2A2axFmzn+HGnYogs7
fXMf1wMj2kC+4YjpduYOIIxTtaZEgbllPCQ7IlaSgR9Vnl+hrWbIhzOK1rWeRX7X
DE9GxMdhxgfHO6SGdxwWpUIZ43AT3Nf39BbhBa2bWFTDfqQ96c2cBEU8IPQR1b8R
R2BNPkMvi7HH7uUNLQ3j1YL0cYcW1eII6IIxYnKjuzIxRBaJyY8hvc2hQ9b1tOSv
YLGCqu3v6/UH/skZA1qB8O4jVKG/bXTC3ZVnMivbXqUkdmXeGjVatVQKodmvv4xN
m0VM4fu58Abj/nemGqF/Qq27LeWJHjF0fnDyjSPE6OP4JVaUUCvAvZ4chxrD0/gZ
uJb3TsiBJS6YJnOJK1EeUALhKOluaxkRdCPWWNSifX/pNe7Wkuf4G3N78EM4bTmp
HYQV058OGWcXJQNprBYaAe4R+4YEq3sfK8jtEbGdNJUpwP/A/aVmujvtwEI7BH7U
1bvwGGXIynJZ0GaHvMdX602+EunmEk1dfZIXN9qrn/31UM3UAcSxw6jU8hKM0jyM
dJZPyJnJOpuvk+EQlXVGOgcVSNO5aElHeuZ3cyxC8iv8V9E+U9E/Aecgj0dmXIF2
8eYyL14tO6KVTY0t4VEabWi7DezrJJc+bBMgb+J0shMJQVXllaogPCqr98a330oF
K7xjeSk4YdXSATQd7q4orqQ9X+9lY+eJLOkjwQGNcrfKrrT+ekvy0IadBfZq0jsY
RjSAMLdbBhf2xNeed2iJwmcvgnIx3Ii0ooG5jHwXRiiEef0Y9YUwCG+eQwEHNxR2
oXhAPmt7421UAn4dsDqhBlRm0x1rLKlQX6pn8Rl5Ktbe73jhU0AWoVSbSRPhcvN2
SHCGzltQdPPsXSmsUJJqVIZsrGkIzlyGhmVH3wqi6H3z/nh7Xm6e/E44EydeiSBv
gDcq5jctxU4LIXk47VRDkC1xtd4WFShL9lub86SghGo0LLRJE0FE2zYTqemHA8qB
XE9eOcYHmWwEDLBSmwEbjgcvE0tawWhGXItsJvB/VC6xHTFCU2oMCYlXo0vK1lpq
UnR7xPIeNIac7EPNYe2/qNL8GsfW/ba04I3YH3+TVgbDP1EPhgDZyD6VX2HpR1UA
nv0Tgv/g3aKdOgGsoPPiJxS9lggDGpLndJ4WbkWgEDBSuzTRseCpxNsF8jUGQUVX
FYvtK/iFz2cvRkoPQAxeLpOUceFaaCVfk/VZdTAe/tM3aIWxgsteUUJ5R9N9UyHs
0tG+J477mY7O1sYzs4xUmVYqmGj9M4WMDmhujxQQq5fnSmoxyR2vAjZW62oapLq/
Cy9hbNYwDxtws0xggXjGIV2O18Ctkt+AXyM6Ab31+4aN0Ll6VNS54Mow8vj2xMQh
gksmVim/eM775qvWYoYDWITQUr345yBlNCjnA1hccadmxI5wjOvpXiws4j4UBF3h
msgxr0wO2eUzb4+baqCD9X7wdmXZX3+oKNt4nUV6+nt/eMOMl/Tvim7+VRXIfq/X
5/Yo0gTQbQ3g5wD6OkznuTinjr8v8OWtQtxGBO5fT+G/NgBTUcTDhpxuavQsfs39
iePHEsKRsHHeBTtU7r3DouzVDe4FJpXAPm2YUgez1IS2KcmWRN/8V1h60CGj+v+z
libx3z3jR/ImZTSRQxXduZzQM8XCeeH3ccGzPhyzzw98Fd9iRGywW+cUdbv0XJpV
DSt+Km1QPxQ0J5BkcOY6iJefW4gY0gBW02rdCY5vXrnl1C6uH4OmgKaySJfB68G4
WG/NxdJU7PR2576EkLLLl4o7bOJersmbaVPKW/GclG8dDXxYd39C8kDfPUb5bYW7
6memHqxfiy+9dm/2ccdyMoMf7QxiHNsqyMuBgZecwThA/dBvlFTMc/az5OSHarHc
5GfzLYhlSzFvowvXqmw1wgH6WtjsdwmZbt33weSLRDFin5TfnCaxMiqFLce6GV8w
jDczjvBiUn5eU49RJuaPXwxZR4aLWCKY9HwEKaxrWA41Whrt7prS/2OTDG0gFGFG
gmj+A1nkbVKlxMiaMcQw6NxXU6g+cRE6hM/P2l14WXQajPnXNrr/r5kotjaUKkuj
obgpf4B9cMav5cHt05OZSmb0v0UQBuldXuBpvFNzFzZX2jHz24cOOkcGV0DKjDc0
o++Hi8gS21eDKR6E2IVeCy/Yud13htv6bgAKAQcd08VM9aS2zuiLMP+rfs8surCb
tUbCBuowh6gOIHodp4CEl2VV3jO/8BocKmXuif1uEjA9NLuOqxAyjrjsBNCmbw0s
3krEMVsXjUlaj7PV5PquNFp36QrinNgeDkJg7DwEtx1WOaiZ1ANrL60wYLpnwEZ/
eOeJ82EcWl5z/NdRRjE9JgsxEYyWLYjtUFH8ySLU1ccuJVl8l2D4/JebGwCa4SFZ
R94+BYHVx5pFoZPIWOG7Ky1I54YsimOwlJF7yP22BCl5dB/+ScWkl1pelD8AmMTF
XyqM469BJoWvdbSnr/QiO1snIPmmN3xTg3R9k8y9vPaUSDbw9/uWXNQhYc4uxuov
cgzb045Fm3exsuSLTAeViUMKbAxKM13jbhWoJmVrbFGH5yVk0SA0M9kQoP5D6Ugf
Rb9hnns1aOHjEnN4T7mng12V6g4+6hOCwM6smMi7TZ5KPeBTxFNSdrfqFgWPU0gk
hBxn2hnzTDl/jcRmAdmttuAYn1TxL77HALoXIMQLXPGHOQ5M8Sq+pYClL03mMaVG
f/p8q5UtoLFI0hXabk0TrE1w+XtvcL71EhylikGO/Oy302NpVIdzoRam4UtRJ2ph
m1A0Tw0y7XGQXk80tJOcr3fa2ifzw2yl3sb6sqzR3arfcvrntElrNPXFsI4qsVGS
zFrtrAhv3YWHl1uP0+a/DGYB9Xe/tE0qk4AMMYYqGSrpm4YAXHHHujQKg7FZaLnZ
h+FfkKq5BnE/FejwGNMe0CqB6cebPWNpa/8f8XY3LhFKPBrBVQrpGgh2NQy360PP
YfAHglaWEi20aO7aJNJ8eQknTxW8t+8+M3aMVzPUeIwXzFKykQt7wJ6QPerMc5oH
ix5OCepNj0MWHJ+zAQLU2t9CCSkueaON8iPEiO1Qin0gzIEB3YKFNopdF2iUEu5n
Vb6TdQIgdjXSlyd30joYO3/14TryDMugQ5c40Zv6ijD09fr6CgmZCLlOF9DY5/vs
G/OZlu+W2uB0rFVop+ZsQrWuyseVSvpXw/xX3CsSW13bfOEycivF4Q4NREF1jT4K
zMhjs0XiMFaMCcmljkfvTdqPhwKwK9YJXPmf8ZCwwhxdi2Aa6xJ8mBC2W+QOO4Z7
jbyq8fo+5Pcm3tAxEkaeqLM/UwQKJjWMnt4TdaFFjo0iBPk7s3gxGivvmqOFS07b
FxTtshXsRlvzY82l1bJWuAWK8/hjixqJ1aSFv8/QrNABp4iUHzD95rNblKUN0K6l
XSJN9xjDOZhHl4IPjQoK4KECASZ+ECAw4cV7EbuCfjWtE7hTs2PhAQRxEhwPPCF3
MJ8ahILlnS3s8Ov5lQYysScy2O3lEfK9vWZscroZMw/rZgb3l3RfNOOMfD5NdZ+g
Po8FOOG/hQRGqfSVWWCLzXVIQTKFl6ByEO8H7hxBg4vk2RqNACpsNe9YePUozbu8
d91am/r0fVvUt0MNrrxcER6C8UsxYHLPL1LDOWiv+PcBrbllbsUFnyCrYKP1Npib
13+YXgtghCTg3MSNOJOvbqQOyI4Zrfyk8MQMbfpIgw/rwD4U3e8qKFiJx1mYQWxn
kZuAdM0dcj3wB+uHP1dIicv82TSv0qD24pVzz4giECXcOTRv2DJ4NLe5F/rTNdqo
9Z34uzPa0u9ZMxX3IIuqyHBA84fNMOsn3oS/vJpFngtTCFvfV4+lrwtvdPSS3mEl
DDc6htcdJFLZ6OaYuL7IakAr74dWijHX9Bi7vSjskMe/gQbV4WH6gK4rHZxVeeDF
4Z1H6qIEZ3zj7UzksUOY0+/k3dwRtAJ37YAWmZZO+4N1SwgdeaIuM1Xc0dj/jgmT
amEfPHW5OYvJj16wWWyB9yJn2o6KIiRKCz2eUf2N2IJnbwgf4ce6jGN/Hk1YjSMu
vMPVoe+buxQPPouXstsBlfcMbD3wtddDcEFgthh9rkcwZWKxXTaLqNPLWwPRZx67
PP17e2Z05jsJaQb03653JkK5w1BJI/BMg7sz9neUxjv5qM0v5a2cToWgZuYrGKi7
7n3apMp5bVFRzWZIkQVoOXuw5ktkLQoxnLEfX6yNhgKcVm3uzCP+XaGHqvBjIZVp
C8DBQ+vRcvK3PMtPBThDJb7KQMR0r2KhjogHvcGT8VVaXTs7Db/RFes10ddSFg78
9KHDymLFaP6aMp6GxjHfZYiZKkRoxgDMdvl34AWp2Jz0ZhkTkPgt/uoLZFhdj/Gy
nsSV2nh/oaKuL++g3o361H+IW/lGFAtUkT923b5SH3v1c0onUdakafDFoqc9UICZ
Et3I5+jBLxAWxm78QeeXsl/tVb0yxPNDApDawWfVgbonXmX8yR3NmofJW6M0MXzJ
8WcMiSWsUldSlftocQ41tZKQfhzYX17HT1S3cAgi3LvM3qAxJqrRIM8QiMmIrVY5
HhElgdsVjHPVwHmYfjaz26Wje7EYvlZ9yn/+c+ey82TWd4TqY6iz8FHU+xbnzd57
uiomzGWVD11QXJH7F/7W+5Fbs1WmUtO0amSLPJ/aZ10buLpueOvGEs363vdYvWK7
kbz9+hEQK4Il2YT9yCYqi3O1W9/YVEcxh5tFCcVLDA4AVYbFo6Rvc8VRd4bpPAz3
Fx54Co3aXJl4+Xs6BJk6pH8SBuW9OaDlsXmgsabjfHVyDmYAq73y0gDjAYCuUxnG
X44UL2QHn9yN/HIzYxpSGten3JDFNl3x0CnW4vPrCMPkXJGaptV6pUo8J+4vUibM
Mpm73Iaau9jvUAjdc8sSUjTAC43XjiiE2bJmge5WyFPIg5+hSpBs22CCmT3vnAJA
AOAH7vuc4sFmT2NmfnUCOErQ/oNPvijj4/9v8DwL7Ptc/sBxo5+25Kl9Ex4jAT2r
ZlQNiK6rucIVU+45p2LgGqE9hJsj4r7woO9flsJrJUHnBJu3dzt6DdNZrm0eWY3i
xO6hbVTYZWyrPuf8EIkoNn4b53ir8iUzOy8PshkT9w/5c2G7XyMOJZnYH8TR7bJu
Ji4rzxk/njOIuxM0DXVQS8zrKI8d0fJTFvWxEHxdEpB0R9w/94tEJsBIvEKO0TI2
on04skCYBIrYaEvPQqF7q8ya98qnsqzZtKjBduHe/U8lOxc0meRsTrIZ29MKdtnR
HTjs1SiqV409bb6hXMvERzb0hChEl0UaN2zVCp7VwkmEXp3yIR3pYJzzry+8krcq
bCzzSgwt7P3RPwcF33cBk2UCVDqO5q4o0rUnrMWQUtYWwkJXQxCUoLVFih9R1S2C
nd517ExN5zx+7osNjUfC73mty4e+H2g/ngoWxzmZjXlHe+bqNcXVTrE2OAkCchYT
gSIf0nlB5h+z/3IZXJP4vd2l1OqUfdPyJ+CQ6FnfATqq+MrKMKxrdEXyQ0IfRtTn
m7LVjWKOEOTd1G90L6vADOyAlKX6hvn/RgMaQDg3HIRalpa48GvYyUQbth1eLOkZ
LmI2yxmaThXUbUfoic1+Kr4u9FksasRoi4DlQdmQIBv6M2378inbbmxgmkRvgMVS
nw3LAt+/xAoLqxb+OGqYJaB9/87Qlfk8cwnACRyxSyh1ghaV2VSyNLHsJ82Uctya
ipmSvcZb+ZEMHfmj8FlEjju4vhH0iY0rJ1JS+IYXhL8nZpj1O/2AUWL+jXSKNrsL
FVP3QdvJ18haPPrtLZWZUdeEnSzg1gVvUAKglb9A1696gXEvNw9eafs0gW3P9EPX
i0/7/QMbGxlks1Bj1oI+uQcplYSorcyXsN5GrYxrqCnIhGBN+GA049sUjiU1cKnG
vnnmqP9kByivG2DYJ3JPdC2yWO+muXbSOEHBqJwBfkOf0KLC7LOptOhSaXQvB8Pb
lhUvEkLhdE97ZjK/mLuWlM5ucHcfYN5L7NsGeVmYuC0yLwBZ07T0txbCpg/LFsEU
zyCq0PuII/XFn+mV44WPxA2DxcZA0N7lljUO6ePGCVqb09RsGfg/1h+swzMuJYNX
PNqJ4IHTmFhvs8QMjcL89oz1GIftbxwzMb+9vclz2lK9s1KvgIS53CtzMoQoG1+v
2AUr5bZMAldgtOiD4MM8xFf97gm299NBFLpHah89JGBz0Uo8A8U2vtCQh89rY/OL
S2MgE+5abtWHL4Oi0TwyrKtuDGYVmglV5sLzx1KQTzlf2j88iJOiOsg48GNqwnrn
I/k/WUNz6NyuaqtUuJo9Yrjr2hKN98eJi8sRzdEzh+chHqvZoWTvd/8djUOi+79P
Qg4JYO6yaIWX2+DKSFQ3Sn/o5o15jr05L+UoWBW5QKWkIvXWsPsUfmR3MwRMDBu9
swArBmHbdwkWMx5rYcgRXiMMoVLSZJZII5lxEHprn6RJXGIur8lMeveWBDMaAdj+
gy9UllsDcGPqYj0c+Un+WWbnvaqb6EWiY/x8VevlgoUrnHfRe1OB1yVOYV31AsbO
5CGOOHy427eJ3kHIEOOcSQnof7aoZ1+vB5JoTNyFUi5ujRTvMxxUAYaZgsWRUMci
FEDwnIttIh0W3XJLjsCWDkUe1v6qBOf8GSiHimFDUYaugszUIwXhcW6UqqN/T25B
GFB9OwTZQshNTsX3Xs8TPNcJy7wrYRAEQJ8niRwfuVxejjH3oRq7MaLLsD8YQxN0
KJQinxBNuxNn+RAX8Lk/cKUfpv4Qw0jqWu9oc4xtVZ5BnkUCwqjKMnmZ+8BA6adi
aldhxAs8CqhUUNtVqPRp81qBT5sy5uVPPKW47cM3XVJFhG75DmXQuJwKieHBIDJH
savsh74WH2vc0JowWVe7ibMUoKYyS3YkudjX9EbBSFi+ThY6W0jK/vlCPocdJqt8
4S6RE7rtgrIrWgCVMs26eetUoM3Eb1yfNKbEktds2SH5awU+eod9bX0hVkcgBH3P
GdXd2eKeQneDVkVpiecLSTz8+dSg4XkFyOGx5+pdf4P5TEllZSsC3+xcJtxoZke3
Qao2sXiyR14mcVVvmiCogdeW+aMjfHoVM1BGq8e6Q0AIJ7ASFAzd2NSXgLLebsfC
D/lYT587+tL8LoYxw4nrW40k5W/eR25GnSjxTYAdVoho/mMUXaud3LZMtqLasxyH
wQMBtVBcwbR+s/fKUu3TOgLXU9h7+a5InRK7cZHbx5+8Ndunjw72/FC43WIc8+1E
qwq+W57RFnd6HkceZSpThmVqlQQ2/NQ8BbuiLzhcOHOs2ks5/eaJv6lg1ByUmObV
Hg9wMCMnB9wuZGOiSpS5r8XlpSrPuTWao/jZssV/yNL3A3W2h/9XPWvnTjN5LA7G
IylNOvYWyBDHcZv9FXj6gnE4xb4TdZ8t38/DLgfE0J/4XDY2LL2IzdNL8W+j8NIZ
Fg+pcSewXLCNTZcyVvlhvjsxspANV5kpHqkhy2rZ+IKBdHrD03yc4obePm4Ki+jb
X3keB+/mVeYY89Fv5qFRX4J50ax7nGPLFoqCvYE0dyCKsnYkyLyXUHxkKEvNXIt4
LfxBN1GSwrrWp39vPS9hks5usP0MW/JatSKQ2XA3wumiFaUuT6P5xScxlzOHNN8Y
8ztA8gWcLoNleviMvSCd+fxmlF6+HSp3TWClIRv3uXzKUmo60kiDCPEqqE1St7h5
Jd3NT+1M7Rsmq79RSqzDCbPew04jmhfD2JFxAN5Zz5nbUZgxHGvKHL9agU1zivns
nOTOOwENq0GjJ/yJvOen8Q0dqAmzPBgWPUxuoVK+JPM3ondurXyqzAdBGDhh9aNI
UAhLfmINZJUOPr1+SDDWe6uMYPeUJFt84g0L9pMIolvsKAUBs2zQS/uO1+mbqgzt
PYRNhBMZd1Qq2r7PF/1cig2sIywZnYcQNSyntH7Q2H58omoEsIb+IvS8he+eZPyo
L3IC8xz8hDVGezTGHgrLDZoOziFvC28IieuldOa8KJHUO82OGiFoM6EAKDa5QGaR
217rx4XSxR3l+3CEtCOWsDIpOpC80os6+U6QPAOxsAMhM4OIkc64q9dlBvGgPfTp
69Ws4jDcXNxTjiK9wsDJE2vWJ+LKGPFz9cloDm1DG1+jC1+DoXgFqbc6j3nWI/DN
AHrfNoCl3nJTPEsuItEys52N+FO81cKYKOda0s9TjjfAZFWF0PXc4w9ljAGKFSk2
6a2rcvCj4qpbv7qU9ro5jvSBq4zF1WvS37SOAhHviLcB+0699ib52zFEwC+66Jz8
/6qqD9VKz+mu5xufIJIHy0A32oggOE1Ws4fytUIwEfnOokoAU4Y4ti2YgyfCL3kg
3t9XXOhgjxP39QnDbgkLibU2mlxcZbaoAjajGhUnVdHsGDyG8QnUxNetXwyIPOi+
OUo1JU3nd1nydQs1ydNRZGlw0ODCd/gaA1TT9jm/hqJqrER0K+nVL/8AApLNzC9W
HacbfHuajJhyL4EmqYnrHbZdfzOvRnPNXEBKbfx14S+HwApMLBQdZMtrKfWqymol
FCqs4t2c1uCGLr+rNnmDrOgDz+fzDBb7HYKVHxctWzbR47Pi7fpidghev6sIxqrD
DoxgG2cIfchqEVd5Y0LYIAelEkgDILrebGxt49Ay9pfwFqzCzFYVvBrPu8TdANrJ
lEy+MuoVUiD4Clo6Z8aGXrEpRQRrq5VieZo9RNuNWeXm2rEIqRspT0W1/JA4/UmR
CbqHRAVyXb7/NfiU5Q4eKG5j+KDOdaVIHdvOXgKMjL+nYzBPq6poWLreY6Wwg0iz
K3q15FMXsTP1i/J4bvkPmispOggs3Gr7ujHZN9bqIevLJvztCjjiKi8PoP1t17KR
YxumJ9z6jBo4pu8ny6vomcuALCaUxfcLg2sjcMB4lUPVamdp1YaYw/XR7/UURl9G
fNNeKny7qlr5b8THXXX2kpYDwq2v8eIgt6kWaAusHHjLOm3HpqM6dRKHMJFZADW0
yfdfSQ4G+H0dhOgzx500bnNmx68jzOo05Ov3hqtHoQ68LHU21LrWzq+mYBpdze2W
/kxwM1zRsUVO6Uu6R54Q2z0E7+enMP77evq9pl+a2Az/zUtKrq+o83M0BeXow3H4
7KZAlCSwR1EoPm6opixiYS80nRol3Qej6cleNe9L6xbSwLQOJCvCE60FInXPY5Jf
7Hutv3O1Z7PJoLaA5KCEjA7E1LUZ7eCGjwg/x91kQ228I3rs6QnWe2GIqrs2KHlW
9CdgO1pRx3z9azOTLwOpdVQmUDcsuuwADFpONFlqtLbYDVrYpEMJa44DqRkM7/Jj
yptPw1xl5nXQMC7KK4lm5lzPseXZJ2Bur1Uu+1wHRPh3kfOuqKLBckcoz1aP/eWI
c9xrDYV1yGe1jqFs+NnRkGpv/KoR0pn/nfEl+U9Q2sollwjFJlEOakMmVbrPggmd
tOxGTKb5B8nUyvIjVSAJe2Ud9ANiesBg+RTJANyS3R3nZlZxn6Z587UkQMCQEmZC
kk65ADn5K4QdZZqmQJYiNBdJ3FrtI9Dcs72sJmyKxwCFtG/KbvmwJpaSQ51xJHY/
QZIBtfq1ADSt3uiuJMwtTB/7yu4GslmG+FcWgf+aDYS4/1tu2h9+gOX9AVpUQA17
h6dqypntO5+onsFs+cFGZoaz9r6/miCRkg0fxs1ihmLkGg2jDK9ZtQrc1/XCV7ES
L7TPagmofZwgxypINAexSY1M3qe4+0+278s10/oMqLJCp+mZB5OmOpxWdKS3RyQk
ln2UtW19C4gx9nxWgNRcxaWXp+DXgy4wrGSzr7CIlq16VMj+aYwL3AwikWHfRVyp
xhBeocpVh7pwH/sdFCryR8NMWefL6GaQI3HO9McOqx139lIVgGJybBuPF5XvRIyy
cbohom18bGDG47ZL7QOrX4/PJcbuMsmhH7TmSFOYi8coW2hxxbOcYs6GicefLj2K
qT2xC+6HLHoIrNYlVlgmOkKBoxMrAalEXiAqUwRT14CaVzXobEvbNzfUCiyYXnoK
z00XTODzdELeZ0FPy+hZm1ybI/z3L7/eeVzZ8ImWDK8dGU6xTElaEVJ0Uf12t/br
sB7iVsv74R4hPJCLl2b50Bx+QVv0AVX0T0OlJIUl9PBVf8TlFaibAlldeqWIOa/F
7BbfW+/bsJ2tIc6ZkAMtZbbAZ43W6n1xRDHV241FcImxA9jRxcnwZzVY1IkRSD2c
xxPWBlcHNppXeG+55qBlQyBMOCLLdFrT7NgFabbH3rmaW+1qDyYocBbLFDrbtMBz
4bJUGPp/8KoK0hppuG2Xr86+amZx500eplRCW/ssmBY7iWQ65xpXLvAA5/n1molX
u4VvMVBarUb20VSrjpVkXuyh5sl65KvL2rDwM0T9zbx/XEONk1c6Sp6HTAu9+0n5
aPax9VCd5OQhCVaJwqmD0aHXAHymLS/QI0zVCg/+eBvu4VFcNw2POoVQMTRYWKR2
2PEMBZq1rmWx9ZQIMpljt62UKQN9dlUYl+Tr/bDCUiQWMbuCEEPH27AHzo3BB6pW
vMt6hrO3Fj+3m/i55ehhNiILf76dINtH7gYk2B3G+SM9vVvne2BHgAbafLnPMpjq
1u4lzri67PCNoCXKQIzZ3kTHrxwTGIV42JOa1p0vsvTX47aVTG3R9fkJlSo2ZZAv
EXpGfs6gJX4coKFMnBXqhd611s/S5hLib8ht9FZi1d+570VjTWpsCn9Bk5CS02bx
msYYKxDREL4Q4dAECtcceKlZreLCPZ88NZKlmicze+pjnLChFVp5JZmfIdDAcwKy
fXe/TtouqlVx47Rd0rzlbmYDZ8AOw+RW/ywo3fTQzFmVEjef+AqHVvfkNOaqHhFE
GEtmt/tQLDzPpslsgQQIRF+H2H1zXbE2lK9U4A51NlkncDdtxLhcpXdxHMnZde9J
CkbYhCHlbQcgrFV4le2ToeTjeBo2q9JmIqSv6Tu3FLun3Vevb86DkeUww06GEYhY
n1dIG2q0Je4g/PSSaapRq9Ewl53Of4ZrueHZdI68tQ5j51RIEf1NRxmIMQ6qY71F
X4lmvF6b41zA/Mt8OTWWznBU0HTnMcEm/HFO/NOF5tZryRuhvmNVCRAOHgJR1scI
Pi46hF0VMXm+bMGqEgBhWOcapiZEn964T8Jl42opBALBQKS7I2Yzx7BBLY6ebNMO
ZYo60cHplATwrm5cKx9tSymygP3V3rMEQ4UQ546Z4ENv2+P87kOapQ7wA4DNZ69A
t/CQNxqs5mQ1S9X6oLLSf0in5amrJUI6D+WSNOZefl2FsVqAjjE3te216MC/K/CR
bwVtkPAoNa5MXRpPOSHRQWxewKm8O/tEUSsica4m9gA3cEZDAC8eYTHvy9VJkYYj
ii+3esA0SVjVhkZrXNRqHaHSmHZDk5vpHK1dSyvj3857KvwQNTHhQTb9RTTJXXD+
WQpjeEj/s6Bu+8AsQb11ABY81N/rSlouQPnPW5NLddXYN8FuUYCkeSsKNW0nBZzh
6wZTNUwdocZLQ53glPmCuLLj5D/51RssDGygWRxSDEvwYlhs7GQO1OfnijfvoygA
CBs1Ol/NQ54X1FVue/SXnOpNmbtqpW4oPQeHxY7XsUBywiFo2KRybcDwe5yR11ll
OhV0xvVbxtuYza7piiBJsuEj8Dt5I0ssiDb/dBLodvY=
`pragma protect end_protected
