-- wasca.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity wasca is
	port (
		altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_cmd   : inout std_logic                     := '0';             -- altera_up_sd_card_avalon_interface_0_conduit_end.b_SD_cmd
		altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat   : inout std_logic                     := '0';             --                                                 .b_SD_dat
		altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat3  : inout std_logic                     := '0';             --                                                 .b_SD_dat3
		altera_up_sd_card_avalon_interface_0_conduit_end_o_SD_clock : out   std_logic;                                        --                                                 .o_SD_clock
		altpll_0_areset_conduit_export                              : in    std_logic                     := '0';             --                          altpll_0_areset_conduit.export
		altpll_0_locked_conduit_export                              : out   std_logic;                                        --                          altpll_0_locked_conduit.export
		altpll_0_phasedone_conduit_export                           : out   std_logic;                                        --                       altpll_0_phasedone_conduit.export
		clk_clk                                                     : in    std_logic                     := '0';             --                                              clk.clk
		clock_116_mhz_clk                                           : out   std_logic;                                        --                                    clock_116_mhz.clk
		external_sdram_controller_wire_addr                         : out   std_logic_vector(12 downto 0);                    --                   external_sdram_controller_wire.addr
		external_sdram_controller_wire_ba                           : out   std_logic_vector(1 downto 0);                     --                                                 .ba
		external_sdram_controller_wire_cas_n                        : out   std_logic;                                        --                                                 .cas_n
		external_sdram_controller_wire_cke                          : out   std_logic;                                        --                                                 .cke
		external_sdram_controller_wire_cs_n                         : out   std_logic;                                        --                                                 .cs_n
		external_sdram_controller_wire_dq                           : inout std_logic_vector(15 downto 0) := (others => '0'); --                                                 .dq
		external_sdram_controller_wire_dqm                          : out   std_logic_vector(1 downto 0);                     --                                                 .dqm
		external_sdram_controller_wire_ras_n                        : out   std_logic;                                        --                                                 .ras_n
		external_sdram_controller_wire_we_n                         : out   std_logic;                                        --                                                 .we_n
		pio_0_external_connection_export                            : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        pio_0_external_connection.export
		reset_reset_n                                               : in    std_logic                     := '0';             --                                            reset.reset_n
		reset_0_reset_n                                             : in    std_logic                     := '0';             --                                          reset_0.reset_n
		sega_saturn_abus_slave_0_abus_address                       : in    std_logic_vector(9 downto 0)  := (others => '0'); --                    sega_saturn_abus_slave_0_abus.address
		sega_saturn_abus_slave_0_abus_chipselect                    : in    std_logic_vector(2 downto 0)  := (others => '0'); --                                                 .chipselect
		sega_saturn_abus_slave_0_abus_read                          : in    std_logic                     := '0';             --                                                 .read
		sega_saturn_abus_slave_0_abus_write                         : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                                 .write
		sega_saturn_abus_slave_0_abus_functioncode                  : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                                 .functioncode
		sega_saturn_abus_slave_0_abus_timing                        : in    std_logic_vector(2 downto 0)  := (others => '0'); --                                                 .timing
		sega_saturn_abus_slave_0_abus_waitrequest                   : out   std_logic;                                        --                                                 .waitrequest
		sega_saturn_abus_slave_0_abus_addressstrobe                 : in    std_logic                     := '0';             --                                                 .addressstrobe
		sega_saturn_abus_slave_0_abus_interrupt                     : out   std_logic;                                        --                                                 .interrupt
		sega_saturn_abus_slave_0_abus_addressdata                   : inout std_logic_vector(15 downto 0) := (others => '0'); --                                                 .addressdata
		sega_saturn_abus_slave_0_abus_direction                     : out   std_logic;                                        --                                                 .direction
		sega_saturn_abus_slave_0_abus_muxing                        : out   std_logic_vector(1 downto 0);                     --                                                 .muxing
		sega_saturn_abus_slave_0_abus_disableout                    : out   std_logic                                         --                                                 .disableout
	);
end entity wasca;

architecture rtl of wasca is
	component Altera_UP_SD_Card_Avalon_Interface is
		port (
			i_avalon_chip_select : in    std_logic                     := 'X';             -- chipselect
			i_avalon_address     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			i_avalon_read        : in    std_logic                     := 'X';             -- read
			i_avalon_write       : in    std_logic                     := 'X';             -- write
			i_avalon_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest : out   std_logic;                                        -- waitrequest
			i_clock              : in    std_logic                     := 'X';             -- clk
			i_reset_n            : in    std_logic                     := 'X';             -- reset_n
			b_SD_cmd             : inout std_logic                     := 'X';             -- export
			b_SD_dat             : inout std_logic                     := 'X';             -- export
			b_SD_dat3            : inout std_logic                     := 'X';             -- export
			o_SD_clock           : out   std_logic                                         -- export
		);
	end component Altera_UP_SD_Card_Avalon_Interface;

	component wasca_altpll_0 is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component wasca_altpll_0;

	component wasca_external_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component wasca_external_sdram_controller;

	component wasca_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component wasca_jtag_uart_0;

	component wasca_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component wasca_nios2_gen2_0;

	component wasca_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component wasca_onchip_memory2_0;

	component wasca_pio_0 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component wasca_pio_0;

	component sega_saturn_abus_slave is
		port (
			clock                : in    std_logic                     := 'X';             -- clk
			abus_address         : in    std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			abus_chipselect      : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- chipselect
			abus_read            : in    std_logic                     := 'X';             -- read
			abus_write           : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- write
			abus_functioncode    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- functioncode
			abus_timing          : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- timing
			abus_waitrequest     : out   std_logic;                                        -- waitrequest
			abus_addressstrobe   : in    std_logic                     := 'X';             -- addressstrobe
			abus_interrupt       : out   std_logic;                                        -- interrupt
			abus_addressdata     : inout std_logic_vector(15 downto 0) := (others => 'X'); -- addressdata
			abus_direction       : out   std_logic;                                        -- direction
			abus_muxing          : out   std_logic_vector(1 downto 0);                     -- muxing
			abus_disable_out     : out   std_logic;                                        -- disableout
			avalon_read          : out   std_logic;                                        -- read
			avalon_write         : out   std_logic;                                        -- write
			avalon_waitrequest   : in    std_logic                     := 'X';             -- waitrequest
			avalon_address       : out   std_logic_vector(27 downto 0);                    -- address
			avalon_readdata      : in    std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avalon_writedata     : out   std_logic_vector(15 downto 0);                    -- writedata
			avalon_readdatavalid : in    std_logic                     := 'X';             -- readdatavalid
			avalon_burstcount    : out   std_logic;                                        -- burstcount
			reset                : in    std_logic                     := 'X'              -- reset
		);
	end component sega_saturn_abus_slave;

	component wasca_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                                      : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                                        : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			sega_saturn_abus_slave_0_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                                     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                                 : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                                        : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                                    : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                                       : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                                 : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                              : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                          : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                                 : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			sega_saturn_abus_slave_0_avalon_master_address                       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			sega_saturn_abus_slave_0_avalon_master_waitrequest                   : out std_logic;                                        -- waitrequest
			sega_saturn_abus_slave_0_avalon_master_burstcount                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			sega_saturn_abus_slave_0_avalon_master_read                          : in  std_logic                     := 'X';             -- read
			sega_saturn_abus_slave_0_avalon_master_readdata                      : out std_logic_vector(15 downto 0);                    -- readdata
			sega_saturn_abus_slave_0_avalon_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			sega_saturn_abus_slave_0_avalon_master_write                         : in  std_logic                     := 'X';             -- write
			sega_saturn_abus_slave_0_avalon_master_writedata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     : out std_logic_vector(7 downto 0);                     -- address
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       : out std_logic;                                        -- write
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        : out std_logic;                                        -- read
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  : out std_logic;                                        -- chipselect
			altpll_0_pll_slave_address                                           : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                             : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                              : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			external_sdram_controller_s1_address                                 : out std_logic_vector(23 downto 0);                    -- address
			external_sdram_controller_s1_write                                   : out std_logic;                                        -- write
			external_sdram_controller_s1_read                                    : out std_logic;                                        -- read
			external_sdram_controller_s1_readdata                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			external_sdram_controller_s1_writedata                               : out std_logic_vector(15 downto 0);                    -- writedata
			external_sdram_controller_s1_byteenable                              : out std_logic_vector(1 downto 0);                     -- byteenable
			external_sdram_controller_s1_readdatavalid                           : in  std_logic                     := 'X';             -- readdatavalid
			external_sdram_controller_s1_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			external_sdram_controller_s1_chipselect                              : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                                : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                                  : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                                   : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                             : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                                 : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                                   : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                                    : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                             : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                          : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_0_s1_write                                            : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                                       : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                                       : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                            : out std_logic;                                        -- clken
			pio_0_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			pio_0_s1_write                                                       : out std_logic;                                        -- write
			pio_0_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                                                  : out std_logic                                         -- chipselect
		);
	end component wasca_mm_interconnect_0;

	component wasca_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component wasca_irq_mapper;

	component wasca_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component wasca_rst_controller;

	component wasca_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component wasca_rst_controller_001;

	signal altpll_0_c0_clk                                                                        : std_logic;                     -- altpll_0:c0 -> [clock_116_mhz_clk, Altera_UP_SD_Card_Avalon_Interface_0:i_clock, external_sdram_controller:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, pio_0:clk, rst_controller:clk, sega_saturn_abus_slave_0:clock]
	signal sega_saturn_abus_slave_0_avalon_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_waitrequest -> sega_saturn_abus_slave_0:avalon_waitrequest
	signal sega_saturn_abus_slave_0_avalon_master_readdata                                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_readdata -> sega_saturn_abus_slave_0:avalon_readdata
	signal sega_saturn_abus_slave_0_avalon_master_read                                            : std_logic;                     -- sega_saturn_abus_slave_0:avalon_read -> mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_read
	signal sega_saturn_abus_slave_0_avalon_master_address                                         : std_logic_vector(27 downto 0); -- sega_saturn_abus_slave_0:avalon_address -> mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_address
	signal sega_saturn_abus_slave_0_avalon_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_readdatavalid -> sega_saturn_abus_slave_0:avalon_readdatavalid
	signal sega_saturn_abus_slave_0_avalon_master_write                                           : std_logic;                     -- sega_saturn_abus_slave_0:avalon_write -> mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_write
	signal sega_saturn_abus_slave_0_avalon_master_writedata                                       : std_logic_vector(15 downto 0); -- sega_saturn_abus_slave_0:avalon_writedata -> mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_writedata
	signal sega_saturn_abus_slave_0_avalon_master_burstcount                                      : std_logic;                     -- sega_saturn_abus_slave_0:avalon_burstcount -> mm_interconnect_0:sega_saturn_abus_slave_0_avalon_master_burstcount
	signal nios2_gen2_0_data_master_readdata                                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                                   : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                                       : std_logic_vector(26 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                                    : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                          : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                         : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                                     : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                                : std_logic_vector(26 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                                   : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_external_sdram_controller_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:external_sdram_controller_s1_chipselect -> external_sdram_controller:az_cs
	signal mm_interconnect_0_external_sdram_controller_s1_readdata                                : std_logic_vector(15 downto 0); -- external_sdram_controller:za_data -> mm_interconnect_0:external_sdram_controller_s1_readdata
	signal mm_interconnect_0_external_sdram_controller_s1_waitrequest                             : std_logic;                     -- external_sdram_controller:za_waitrequest -> mm_interconnect_0:external_sdram_controller_s1_waitrequest
	signal mm_interconnect_0_external_sdram_controller_s1_address                                 : std_logic_vector(23 downto 0); -- mm_interconnect_0:external_sdram_controller_s1_address -> external_sdram_controller:az_addr
	signal mm_interconnect_0_external_sdram_controller_s1_read                                    : std_logic;                     -- mm_interconnect_0:external_sdram_controller_s1_read -> mm_interconnect_0_external_sdram_controller_s1_read:in
	signal mm_interconnect_0_external_sdram_controller_s1_byteenable                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:external_sdram_controller_s1_byteenable -> mm_interconnect_0_external_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_external_sdram_controller_s1_readdatavalid                           : std_logic;                     -- external_sdram_controller:za_valid -> mm_interconnect_0:external_sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_external_sdram_controller_s1_write                                   : std_logic;                     -- mm_interconnect_0:external_sdram_controller_s1_write -> mm_interconnect_0_external_sdram_controller_s1_write:in
	signal mm_interconnect_0_external_sdram_controller_s1_writedata                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:external_sdram_controller_s1_writedata -> external_sdram_controller:az_data
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                                : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                             : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                                    : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                                         : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                                          : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                             : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                               : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                            : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                                   : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                                  : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect  : std_logic;                     -- mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata    : std_logic_vector(31 downto 0); -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest : std_logic;                     -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address     : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read        : std_logic;                     -- mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write       : std_logic;                     -- mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	signal mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                                          : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                                              : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                                             : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_pio_0_s1_chipselect                                                  : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                                                    : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                                                       : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal irq_mapper_receiver0_irq                                                               : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                                         : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:sega_saturn_abus_slave_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sega_saturn_abus_slave_0:reset]
	signal rst_controller_reset_out_reset_req                                                     : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                                                 : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset                                                     : std_logic;                     -- rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal mm_interconnect_0_external_sdram_controller_s1_read_ports_inv                          : std_logic;                     -- mm_interconnect_0_external_sdram_controller_s1_read:inv -> external_sdram_controller:az_rd_n
	signal mm_interconnect_0_external_sdram_controller_s1_byteenable_ports_inv                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0_external_sdram_controller_s1_byteenable:inv -> external_sdram_controller:az_be_n
	signal mm_interconnect_0_external_sdram_controller_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_external_sdram_controller_s1_write:inv -> external_sdram_controller:az_wr_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv                         : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                                             : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, external_sdram_controller:reset_n, jtag_uart_0:rst_n, nios2_gen2_0:reset_n, pio_0:reset_n]

begin

	altera_up_sd_card_avalon_interface_0 : component Altera_UP_SD_Card_Avalon_Interface
		port map (
			i_avalon_chip_select => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  -- avalon_sdcard_slave.chipselect
			i_avalon_address     => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     --                    .address
			i_avalon_read        => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        --                    .read
			i_avalon_write       => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       --                    .write
			i_avalon_byteenable  => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  --                    .byteenable
			i_avalon_writedata   => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   --                    .writedata
			o_avalon_readdata    => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    --                    .readdata
			o_avalon_waitrequest => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest, --                    .waitrequest
			i_clock              => altpll_0_c0_clk,                                                                        --                 clk.clk
			i_reset_n            => rst_controller_reset_out_reset_ports_inv,                                               --               reset.reset_n
			b_SD_cmd             => altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_cmd,                              --         conduit_end.export
			b_SD_dat             => altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat,                              --                    .export
			b_SD_dat3            => altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat3,                             --                    .export
			o_SD_clock           => altera_up_sd_card_avalon_interface_0_conduit_end_o_SD_clock                             --                    .export
		);

	altpll_0 : component wasca_altpll_0
		port map (
			clk       => clk_clk,                                        --       inclk_interface.clk
			reset     => rst_controller_001_reset_out_reset,             -- inclk_interface_reset.reset
			read      => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write     => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address   => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata  => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0        => altpll_0_c0_clk,                                --                    c0.clk
			areset    => altpll_0_areset_conduit_export,                 --        areset_conduit.export
			locked    => altpll_0_locked_conduit_export,                 --        locked_conduit.export
			phasedone => altpll_0_phasedone_conduit_export               --     phasedone_conduit.export
		);

	external_sdram_controller : component wasca_external_sdram_controller
		port map (
			clk            => altpll_0_c0_clk,                                                     --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                            -- reset.reset_n
			az_addr        => mm_interconnect_0_external_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_external_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_external_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_external_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_external_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_external_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_external_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_external_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_external_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => external_sdram_controller_wire_addr,                                 --  wire.export
			zs_ba          => external_sdram_controller_wire_ba,                                   --      .export
			zs_cas_n       => external_sdram_controller_wire_cas_n,                                --      .export
			zs_cke         => external_sdram_controller_wire_cke,                                  --      .export
			zs_cs_n        => external_sdram_controller_wire_cs_n,                                 --      .export
			zs_dq          => external_sdram_controller_wire_dq,                                   --      .export
			zs_dqm         => external_sdram_controller_wire_dqm,                                  --      .export
			zs_ras_n       => external_sdram_controller_wire_ras_n,                                --      .export
			zs_we_n        => external_sdram_controller_wire_we_n                                  --      .export
		);

	jtag_uart_0 : component wasca_jtag_uart_0
		port map (
			clk            => altpll_0_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component wasca_nios2_gen2_0
		port map (
			clk                                 => altpll_0_c0_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component wasca_onchip_memory2_0
		port map (
			clk        => altpll_0_c0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                --       .reset_req
		);

	pio_0 : component wasca_pio_0
		port map (
			clk        => altpll_0_c0_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			bidir_port => pio_0_external_connection_export            -- external_connection.export
		);

	sega_saturn_abus_slave_0 : component sega_saturn_abus_slave
		port map (
			clock                => altpll_0_c0_clk,                                      --         clock.clk
			abus_address         => sega_saturn_abus_slave_0_abus_address,                --          abus.address
			abus_chipselect      => sega_saturn_abus_slave_0_abus_chipselect,             --              .chipselect
			abus_read            => sega_saturn_abus_slave_0_abus_read,                   --              .read
			abus_write           => sega_saturn_abus_slave_0_abus_write,                  --              .write
			abus_functioncode    => sega_saturn_abus_slave_0_abus_functioncode,           --              .functioncode
			abus_timing          => sega_saturn_abus_slave_0_abus_timing,                 --              .timing
			abus_waitrequest     => sega_saturn_abus_slave_0_abus_waitrequest,            --              .waitrequest
			abus_addressstrobe   => sega_saturn_abus_slave_0_abus_addressstrobe,          --              .addressstrobe
			abus_interrupt       => sega_saturn_abus_slave_0_abus_interrupt,              --              .interrupt
			abus_addressdata     => sega_saturn_abus_slave_0_abus_addressdata,            --              .addressdata
			abus_direction       => sega_saturn_abus_slave_0_abus_direction,              --              .direction
			abus_muxing          => sega_saturn_abus_slave_0_abus_muxing,                 --              .muxing
			abus_disable_out     => sega_saturn_abus_slave_0_abus_disableout,             --              .disableout
			avalon_read          => sega_saturn_abus_slave_0_avalon_master_read,          -- avalon_master.read
			avalon_write         => sega_saturn_abus_slave_0_avalon_master_write,         --              .write
			avalon_waitrequest   => sega_saturn_abus_slave_0_avalon_master_waitrequest,   --              .waitrequest
			avalon_address       => sega_saturn_abus_slave_0_avalon_master_address,       --              .address
			avalon_readdata      => sega_saturn_abus_slave_0_avalon_master_readdata,      --              .readdata
			avalon_writedata     => sega_saturn_abus_slave_0_avalon_master_writedata,     --              .writedata
			avalon_readdatavalid => sega_saturn_abus_slave_0_avalon_master_readdatavalid, --              .readdatavalid
			avalon_burstcount    => sega_saturn_abus_slave_0_avalon_master_burstcount,    --              .burstcount
			reset                => rst_controller_reset_out_reset                        --         reset.reset
		);

	mm_interconnect_0 : component wasca_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                                      => altpll_0_c0_clk,                                                                        --                                              altpll_0_c0.clk
			clk_0_clk_clk                                                        => clk_clk,                                                                                --                                                clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset           => rst_controller_001_reset_out_reset,                                                     --     altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			sega_saturn_abus_slave_0_reset_reset_bridge_in_reset_reset           => rst_controller_reset_out_reset,                                                         --     sega_saturn_abus_slave_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                                     => nios2_gen2_0_data_master_address,                                                       --                                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                                 => nios2_gen2_0_data_master_waitrequest,                                                   --                                                         .waitrequest
			nios2_gen2_0_data_master_byteenable                                  => nios2_gen2_0_data_master_byteenable,                                                    --                                                         .byteenable
			nios2_gen2_0_data_master_read                                        => nios2_gen2_0_data_master_read,                                                          --                                                         .read
			nios2_gen2_0_data_master_readdata                                    => nios2_gen2_0_data_master_readdata,                                                      --                                                         .readdata
			nios2_gen2_0_data_master_write                                       => nios2_gen2_0_data_master_write,                                                         --                                                         .write
			nios2_gen2_0_data_master_writedata                                   => nios2_gen2_0_data_master_writedata,                                                     --                                                         .writedata
			nios2_gen2_0_data_master_debugaccess                                 => nios2_gen2_0_data_master_debugaccess,                                                   --                                                         .debugaccess
			nios2_gen2_0_instruction_master_address                              => nios2_gen2_0_instruction_master_address,                                                --                          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                          => nios2_gen2_0_instruction_master_waitrequest,                                            --                                                         .waitrequest
			nios2_gen2_0_instruction_master_read                                 => nios2_gen2_0_instruction_master_read,                                                   --                                                         .read
			nios2_gen2_0_instruction_master_readdata                             => nios2_gen2_0_instruction_master_readdata,                                               --                                                         .readdata
			sega_saturn_abus_slave_0_avalon_master_address                       => sega_saturn_abus_slave_0_avalon_master_address,                                         --                   sega_saturn_abus_slave_0_avalon_master.address
			sega_saturn_abus_slave_0_avalon_master_waitrequest                   => sega_saturn_abus_slave_0_avalon_master_waitrequest,                                     --                                                         .waitrequest
			sega_saturn_abus_slave_0_avalon_master_burstcount(0)                 => sega_saturn_abus_slave_0_avalon_master_burstcount,                                      --                                                         .burstcount
			sega_saturn_abus_slave_0_avalon_master_read                          => sega_saturn_abus_slave_0_avalon_master_read,                                            --                                                         .read
			sega_saturn_abus_slave_0_avalon_master_readdata                      => sega_saturn_abus_slave_0_avalon_master_readdata,                                        --                                                         .readdata
			sega_saturn_abus_slave_0_avalon_master_readdatavalid                 => sega_saturn_abus_slave_0_avalon_master_readdatavalid,                                   --                                                         .readdatavalid
			sega_saturn_abus_slave_0_avalon_master_write                         => sega_saturn_abus_slave_0_avalon_master_write,                                           --                                                         .write
			sega_saturn_abus_slave_0_avalon_master_writedata                     => sega_saturn_abus_slave_0_avalon_master_writedata,                                       --                                                         .writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       --                                                         .write
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        --                                                         .read
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    --                                                         .readdata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   --                                                         .writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  --                                                         .byteenable
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest, --                                                         .waitrequest
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  => mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  --                                                         .chipselect
			altpll_0_pll_slave_address                                           => mm_interconnect_0_altpll_0_pll_slave_address,                                           --                                       altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                             => mm_interconnect_0_altpll_0_pll_slave_write,                                             --                                                         .write
			altpll_0_pll_slave_read                                              => mm_interconnect_0_altpll_0_pll_slave_read,                                              --                                                         .read
			altpll_0_pll_slave_readdata                                          => mm_interconnect_0_altpll_0_pll_slave_readdata,                                          --                                                         .readdata
			altpll_0_pll_slave_writedata                                         => mm_interconnect_0_altpll_0_pll_slave_writedata,                                         --                                                         .writedata
			external_sdram_controller_s1_address                                 => mm_interconnect_0_external_sdram_controller_s1_address,                                 --                             external_sdram_controller_s1.address
			external_sdram_controller_s1_write                                   => mm_interconnect_0_external_sdram_controller_s1_write,                                   --                                                         .write
			external_sdram_controller_s1_read                                    => mm_interconnect_0_external_sdram_controller_s1_read,                                    --                                                         .read
			external_sdram_controller_s1_readdata                                => mm_interconnect_0_external_sdram_controller_s1_readdata,                                --                                                         .readdata
			external_sdram_controller_s1_writedata                               => mm_interconnect_0_external_sdram_controller_s1_writedata,                               --                                                         .writedata
			external_sdram_controller_s1_byteenable                              => mm_interconnect_0_external_sdram_controller_s1_byteenable,                              --                                                         .byteenable
			external_sdram_controller_s1_readdatavalid                           => mm_interconnect_0_external_sdram_controller_s1_readdatavalid,                           --                                                         .readdatavalid
			external_sdram_controller_s1_waitrequest                             => mm_interconnect_0_external_sdram_controller_s1_waitrequest,                             --                                                         .waitrequest
			external_sdram_controller_s1_chipselect                              => mm_interconnect_0_external_sdram_controller_s1_chipselect,                              --                                                         .chipselect
			jtag_uart_0_avalon_jtag_slave_address                                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                                --                            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                                  --                                                         .write
			jtag_uart_0_avalon_jtag_slave_read                                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                                   --                                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata                               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                               --                                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,                              --                                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,                            --                                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,                             --                                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address                                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                                 --                             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                                   --                                                         .write
			nios2_gen2_0_debug_mem_slave_read                                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                                    --                                                         .read
			nios2_gen2_0_debug_mem_slave_readdata                                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                                --                                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata                               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,                               --                                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,                              --                                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,                             --                                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,                             --                                                         .debugaccess
			onchip_memory2_0_s1_address                                          => mm_interconnect_0_onchip_memory2_0_s1_address,                                          --                                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                            => mm_interconnect_0_onchip_memory2_0_s1_write,                                            --                                                         .write
			onchip_memory2_0_s1_readdata                                         => mm_interconnect_0_onchip_memory2_0_s1_readdata,                                         --                                                         .readdata
			onchip_memory2_0_s1_writedata                                        => mm_interconnect_0_onchip_memory2_0_s1_writedata,                                        --                                                         .writedata
			onchip_memory2_0_s1_byteenable                                       => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                                       --                                                         .byteenable
			onchip_memory2_0_s1_chipselect                                       => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                                       --                                                         .chipselect
			onchip_memory2_0_s1_clken                                            => mm_interconnect_0_onchip_memory2_0_s1_clken,                                            --                                                         .clken
			pio_0_s1_address                                                     => mm_interconnect_0_pio_0_s1_address,                                                     --                                                 pio_0_s1.address
			pio_0_s1_write                                                       => mm_interconnect_0_pio_0_s1_write,                                                       --                                                         .write
			pio_0_s1_readdata                                                    => mm_interconnect_0_pio_0_s1_readdata,                                                    --                                                         .readdata
			pio_0_s1_writedata                                                   => mm_interconnect_0_pio_0_s1_writedata,                                                   --                                                         .writedata
			pio_0_s1_chipselect                                                  => mm_interconnect_0_pio_0_s1_chipselect                                                   --                                                         .chipselect
		);

	irq_mapper : component wasca_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component wasca_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component wasca_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_external_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_external_sdram_controller_s1_read;

	mm_interconnect_0_external_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_external_sdram_controller_s1_byteenable;

	mm_interconnect_0_external_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_external_sdram_controller_s1_write;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	clock_116_mhz_clk <= altpll_0_c0_clk;

end architecture rtl; -- of wasca
