// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n9D7vbfnOraXKM47OpBEmHL9URfeZ4Q8HSuhBpoVnqvmdtpM93b2crtaph25yjfj
q9QhyAphCe/r6+zGFfml7jEzGrD5l6J1ODCcWjDGG1AyGyy6FJt5vt6TeZ5BpiY3
67Yg3g7UExZDQaM+oqjVQrgL3Btk02Mubjwn+FJk8sg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
4oDJMvZ31gMud3PRAuXlJTB8+iE5JvrpHOe90Fb2CqP1WWAlc+K/bPVxS4edZObb
w72zBkgU+1+jU099ROqod8cR73AHCqFGtTYEC3gmO+6j1cBDh+YFk+Pbs7kZLgCb
PLxT4WkSLjwByErxjYrfl1wE4Hn863E+3+ieSpD9fWlP4Q3yQiqKnre7jh5+ML4H
Uro4+tCBlnRyRPQ15IEXjq6NwoK5kpJSw4PriILpHOFbQ883wlI8BM3kVS/7Tlcx
uHZ0kxrCVoQ5rHEqyjhcrqHcs9ELYr7v+gS8Sj1ShswMEFpAxBYhQq8gTK5VOO57
yWTM0ILZG4H51ieqn2cgr32r/9bOzidLBAszXuHiQHY3m5Kv/VyR/R2VvWKJIjOs
ufFzS0b2lCksgTij1vZ1JC1sG1eO4lkrNTIGcB5qFJgmjr8NK1OA3aVRg2+D8l/U
1OrfoWvLSXRPEL9HbbcZVhe7brcXG6JdzqvO4JOktXGCzPVDVNA57Dxd/yYf6UNC
/ijVAEz1wG/jkWvqj3OLtlVOSXQRb9v7LdyQOxI1XMws1q7SKS3ypHd36yk4p7hg
oXtSMfYXcMD7j0N78XzJzxhMiLYuPoWDNEku3YBEprgVYT7nrwN5XUL144hlNRwF
o6uAY36/db7ymrDtL3TUZC9bTbJxwrsT2b1jDMGDcOa6BFetbkZoDTfu1qeIjDEK
PIxYLDq0B3V9v2P/bkYAdohEvOEdc+O1qRMtVQZKKGbhaZyORCZANJNy55TnsE4D
Rm5dvwoSVRSvJjrKEjH0bRgIzktZCR7wkxhhUqXuJSxyU/d4kqM6dhs5vkvgIaFd
MseJgty/8w9gZbOlungbRMAzI2uZ57RQxeDNxM/zCDFVJ9fSx5FRe4E6acE05NLd
q1Id8s+Lv5StLeqnmkI0JewOjjuFCcsmE3I0pXxp1AUItMFRyBFZyc4YRucyfBUW
fzZFUnAclqgd86P5SfajInqMcT1xITKq84GPdT19KPS55vPdepbVojGPe+Kvg18q
+Kvi03NsdVNdr1qjNcIJmXMxaRPJwdlaTQHOM6iE2tFkwS+m+i3ZJziEzdvW0sNh
8npkfeWPnJMZbt98wa1JjZ2jtSAjTOy+oAJlea9HPVct/sTx1vM/Nto1C9xDg3O7
wwR06c2zj6egooAuGBOdEOAeHgZd5wdJnd2xZLvHhW4/7wDafj39ex+BgGtsMn5j
UAu5bi7M4pZvcXqr1QyLT9xF4GeUW4AMUvCKCFVBpFose5fW/kIHcZJ0ASOdswdP
SMN/fowrFuxglymRykJ+fehtlUXcSdYOJ54h3li0U9EL+GMXklnhx6fUWgB6FG7G
h5EFMmMaWgGL7PQdDajOLgO/d8MYwe0WmtjbdyCcrv3nUfQrLRuT3n+0XgRQ2qrF
6iCQbw6sUUiNynJ0//gN8Ho6Ozq7yYqAX+Wh4+dZeB8+S2bTqMF/w5q/x68kiJdW
4u7dTfVTCFbDRyH3cEyRxXuS4CgZZPirNDgRT+Cq5WGjwJ1LKQxFobrUfBl7ah5D
6yYX+iyh6Y5PFXFfY/vGlRWAn+DOGGb/i7I607AG8m62cNRIj36iCARpTbp8ASN+
+0PB2DUJVYoEDVtswXldKqu6M7IfWVsCHIdVQqzV0gB/EmKH+IIRqufgDyPwhF16
BTn1n2Bp3p2WQs0HIT9z9hspsU29hLbRVvzU8wRoX8rhZb8sZ3WKRKRTsumki+LX
STraQuLlKmJE4eEVybQoVR1QzbUwKN9iDt7k8JzJMU6CyzkbOyJxa3gQz7EeGVNs
cHJrWZtD8auRj0bMd/j8shm4o0Tq7ulJveYjHO7spu8vytBOELJC6XjT9dG3U6gR
pdrEzg7uAMbkYJCcixRQWo1LqTUrmT2RbxaeMQGYmR7N1dnN1vjJGgvQ8ypSY2r3
cvYPRcRWpEvNPHUrXAQbMM3YgjU4xbAwVWi4Kj2q2NhWqEL6gFoKQN+CpvJYJjCZ
k2pXX5ytjniCtM7LicUQQWZJsYWKm/z3NmSpwtjNh05P1FLxckgPF5YTZfVoo9xb
VK7loYGJlpoVSGRgbGsnrapdVelCdhb2lym/6mhZ6KmsCqBT3voEJbfXo4uBqQ8R
1Bi3md1rg6DDj0MFos+bnDL0/mok4nXAi0N2Ko/DPuUZ8I1nLzQCL5T3xUN6C1kV
T8xaGgmJENQP/G9L/Bg64avQwZyIQBCYibOJsGos/WZ92cYIk/fnu63+QmGwzwIJ
e/+2vsh3x8Sg+GryTV4DAYRXZwYyArwyNMfaTXJm6ub0deaGpEkUfm1MNLo9sx32
AqgzUn7EVRrnRyp0ZhKJepSSB4w1Hm6HfV/fHYU9j79wCwWJq5j5U/ya5Z/XAnis
Ni3KSWBlFsIFuRs2fpp7ZkY59xbNWEKG2YWbKJMCgA2FzPU2PBEZ8EWzMTnMGN4v
EqVovw6OwRg/2YKZ3JgA17iDg06wG+vRGcOaX3UtZ/CTJag3TfMAP/Ht6Y3fpO4K
xaEzncZhZzPU14bfZUCOtluemg4FGAwbTrbUPUrT0b2mfEOTP0HIQpTCGVl4H/br
YrMQoSrv3n2rq2QVirHI2tI9sugQENnKrCwBGVZQMI+r6uUjzkoOfic6EsIBD6Gl
0tLPWUNu2VGe89fh6riz+jDJCs01JrHsKQToIR4QVnhcw1Nw20Hx5zLi4Uh3T+Yw
ZV5nhfAFv33LONrcncifkeH42D5t41fDzNLoxi0cjfCsZgfzkNpPt4xS4nQHhtYF
miLKTXmLQeGaLfKJF5nWeihESMh2qTMGNRjl/r5B59WUY9vIE/M69YklyK/G53ad
CuOEcyTxrBehFLS4B3mk9w/ZUarxHMxTgO5rfABcB4ibAHCGuQvCqbCZmXxgcZ7V
woBEoVr9p9TxCNIQoBAlmss/XkscPVZ14EXVpLJ6l/DFI53XMM2IkbhJ13S7lYXZ
yvaF/VXUqdvlXWE42KCxSpW4aps5NhXuUn4wBn6jmDXARQd5vJcycdJMCwFLRjxt
yKiQgUrYqSsESyOlTZPQJ0kuhwlePDbhKyOpe689DRLJAPNvzYekNmTDajpqR/8h
lY03Hsp38k78ZGNULMhyzGtfxU7+asHOsl9mCcoF9tTf+A9BNT94fgwEgMEEO//A
VcjJabnVFOHnmDvgz3R3fg4jkx+w8OwMb73k90LlhGpCHSPQagGLAaQfXK316YVM
y5tsdT+dUNcrnotp23iVs/VAmwX3SrhJsEWyYN/JhqUExAW5tWoUgD4fRncS0nbZ
Fm/m4K7Nf6vFPb1hyDOMj6l0GRNxQuoZM3C0BkDtErBQCF+/GLk8y6VksQgJleEP
a5pA929iJuMiCFvmDRQWvTMcjlaIWtb38/bjrZEMfn/8SOZKYvwSSeAHW9cngMKK
Y14L1kMRteZNuuvK1FhkbGj+9UDUWvTyuOgArEiBWf+7SzI745bL6QDwqT/sgzDd
ZKwnI6/r8V6+P4Li4h9BK3fQF53W1/L6bUPC1i8Z167n/tKRkvSIhtCLM9qDRazt
9SJauozUX2J+WUDNMAiYUc6SIlJBWpOvwPpJwms5IraguC/mbxBKgGDGzFoHi5/j
shVGPC9ZSK5XH9CKseVv45rZKaVJ29jmSs+VyEtMuVve5hIHk2NUSV3VpAtatYgK
R8I/ivC14oDJLYlyvfUCMAv2pBqyQlT9AGzkKIN0+B8xwdQzpztObwvWXS3kHqX6
4NvWG42xcnf/eAwyEMRTDPWVxAtx5Mrw8NIfM5FkdEbwXfjlZgRK4siEYGCSdQqc
hJbT9taFNIhGG0K/92Sp1WiPTC/AdNdt2nKgQXVpIYvaxyXPbSZ6aBv61W0pvgCn
G/6XViWQAWA3EEf11FdgY7ynDeB+0UL1r79YGxxAjjyKgQ8CW/Jlj6aNLxIdH7/w
fptA4XhqQmrao+9PbI3ftpWyOi5YZIYTouqphjyE9S9Oy0lSTDeWFeUyu99fgL88
M0jFaFfyIhd6bFVb+OQsWPqR5lu0reMxCnzKwym+VSowO3CIB65/CxgneojU6cle
Y5mh/42c1b7humB6p7s+AiVQS7unz41DiApsBWNFfCLag42FMcRgc7nXsvscrjdN
I/T7HxRjTWglFXmYI8Z9/W8Ls4gCydKZPDqXmGxLM56tBe/rrHYPP67qL1DORcXS
4JXfJqQgAkPOz97KpvlzevMr4dX0mTGZjdNrFOje6OwPX9rH8iVaULbFMI0xVWMu
8zfypiHkuSaCmBMAcPI5QqxFnMOkf8UrvPvMM5I5Ca1pdtqYwPuFIJiWJEzlE/Gg
Cce+ArRoGIVBDlNyTYhE2ZbGNSTSygsl3XG0CzSQF76XfPeOzHXh1MMwyAoBNloK
YshFzugio7dr4MSbn5aZZFGafP1Q1+p5IpqsS88BJssysbM+pWbmK5ueXGsYJUyr
St70HuXXrSDIN6b5FxrmIX3WmsGVvX3BYXXZD4y1ZE8j98qYjtbReWl/oXvFEi05
R6erp7ylJfwgcF3FDaJ7I/sVVO9z0WGQRk9n2Ud83XlNq59o8er9QLw9/m5gP/nS
usrYcN3rPfBeGR3T+TO+tz3SjWMoI2XmZpijXVGlv+bb2GhsfryY4l8cvDXGJQtn
EF1v5dJzmG3PU52z5fcMtHcUcFQNj0D6xBmKgpUqV/U79bUao6dez3Ua+Qaixkw5
WkpxGpKt4C8XNzoA6Pr3nKdDP18KFFPNanHjTm843HVhjyDAjfpRShZA4L55eIgt
aBx/1uq11ri8bbN/TOFKiijfaTASXsyNMWGnVcM0MUguctocmmGNx0fs9eBL+1h0
0U4DGyDFPA3vJn/N2Auc9WSY4WJlpet3cCcKI2sCwi1cexC+qsbhl6DybufsHztO
7s/4N6oJPtayzWNcV2Gj7+T8Wvscv9WHlL/MbGyg03t3u0GRiKsBhKMo6U5j96Cu
Dm4B2TxEVkyKd8X43EYYT3EYDeo8s/eUu7DbwNmNQwoaSr0dzHaN1E+FVTXO3xxw
4cdxtNB0Iu5NBGTADUV14hSPZ+tN7geh1wkn9+zn3CU94ipxycArFfO38JXP+uLK
OMxeg3s1umQY6liJu15NNfNlFuy3+HtXUYKkjZTLt5gXTNYUXzyhwkj2SEzZ9ssk
NV72dgCDTPVTwzUsPKscYUJXEX1nyxmSMFIgKvxEBvmv4LSQ+wghYOJSApMG7Hja
N2YsslRs0ZGvzV5j2ElAzqJ6KklYfM2GKGJGVhpgwd7hlC77ZkWD/HORWVzmH40j
pOZovJ7+X8iBnju2T5vTbi/ucaNZvwFlT5ES7643/cYdNpUOxr553UcKSqPPyp0c
1/cJoFu7wQCotVYAbbEZ5KE8ATLIIDxBrIV/GNWfAnlDaA9dCyojeOnh9dDwOCdG
MOfsnWK6Jy7VQEiJ0FNkzNxBumHrROI5YP2ATZKsWZ34utXaprGtQvemmCAZMXoi
raR+/5bSzfWVC/yIaC2wXkOIPczYQ6j/Ha8DtJnUhRAhFy8Whxmb4YPUeAcz6++b
3vb57a1mK53SIxK/iF2SeRB9VsfcUSW/hJyiKZPG5H9weLaO3R5PYj/PXskHuSKX
wy7Xwt418WGGfjdEVZ91qedfA1NJZsgZoHBzD2+sf1rMcL+Tspy1TkmamiH36nt0
/4D4T3V8ckk1jme3mjN5i5Rv22GHJ8c1arkk5vNabmwIKPCwvanDFfLLrssTCzhU
sx9y2p1uViAl7ZrSRLhJ0ESC/Bv7Fze5xoH1No9649dQNWhg6+m/1E/Qj7rIGqVx
rkz5uJsbMrygMsLb4llEWGtrSMYRJxRgYE0S4jScjmcfifaS4Cvq5QW1srIPGmMR
HIrqRXqeBsSzQ9eFeFV2M9iSg5SRRUvbF4rsdJl/wdWJ3MPL7ZdhFkDwVO8TuR4a
jWUC10uulIycEc7xy1IjusduX9LV0gVmPAs9qEpu1AchMoOH/+pEpARoT5UWfWGW
3ZYOUfWgKarHh9EvQMc/CliR5U+C3ioXnoAgOr3YQD/f+fNayQL1PdtoTrc5OXVN
WBXWIRlRJ64l4e9+IChGaJMZRO2m+Yjp41NJsFxCEO9biQ2VUKAAEAwHRNglXwNY
rNkuXlpo06O64FJiHDWl8DPb5J6PyZDqr2a3sGfjx0l8IiVtvttapk3Zgtu2Cv79
HxIWr8pzu/vnUg4cq3VMlmBbUZGjTqKc+cocwzFvGpnf4++FVeFZzLX/CCg7/2Kk
MA63ICZoHtgvu2Ahai4EQybyjjpdwc72PA+Lr5Qgc+ekf8TB8UMajARd3PNmFVkv
8Gx2DyP5yz5ISBrDYqtF/uYrrA11cqwL+43ihG1cUUJI9SaM0hDyThreJ/h9NQi2
h5iFTqe/XQ8RvPpda0iXA9iCzvm1pcIT/iTf2XQtqcLaqbtRMLvTl9BWSrhhvNe8
pR8uC46biMxw2T3cSgbkZrlHe5byN9eqcwOgDqqowxEin6qpeKOmUoH+rSkmsHhG
ynAnPnMck/h7RGFS0blN1ho4T4RAEjTxVPT6pvlgskBL5vqzXMhiYum7++BF1usx
7Q2IzoAA0kNf1+VJZpNwFU9wmyUNxU6lFCV5DcXrh6tVBd5aWqWeKvjwsNNColbQ
osPQ8ZDTPjPcHgCzImiA9LR2glC/2nFA9CuYRM5DeHwAnK9jhF0wdUXU+bIMXIyG
ttb/0nso0vw6RZHotQbe1K1lUil6YC9JfQW8JnVm6yob9xhWbZVePVA6o3aE30dB
XfPqmKCnUdL9Nthwi+4ctQHhvaHvFa1GyyKFE/ip5NbvBDzFzzkSPfqdhWztj0/R
jwNif3K354ATCwpwX0iNjhm2WaZmrCrukD49lEN2/DArZ8K8GbEksDzvU8CKwDT+
FT6KGxOHWFGLSO2JJSqWjlzd2bvXkL9WFxu2I92xBFkZQ8vMjk4DXLU8aCFxwI8x
eT6xphs4jY4YG30mQR9uzu0NhjTmvUuKwC/0zRar25xl1g/pXcxAOtJKH+nSse++
SFRuQWVW0I7N+73qvBH5Ws0udPm21lVdEE3PZZR0JF1Uz3WIKRRdF3EG9c98yLbN
aKHcqSoLdQnvbTr+wLpmCq1cPjx/O65oYUh3plc/nJxrxk3EDwTy+PxrqMhRDNYY
1qrnyEvKIIFhHmtJtThWt/RlPbQQlojOlGW4WiYOBIihaShcjEipzuQcSgOg0fUo
zki8oWTHrwospRziVES9Lsx3F0ZnifTSDZPG4oFfhhRGfpci1V2dYWRWnHi+N5du
6Ox1joPa8MOMhCdUvWIvK3VnF3RMNLpdLKahJ82a2LLaZgCsba/sqQnXbTinEUzv
gahDs6ejJ/0CeGnu14AVV0GfVY1FLM59zpaSOFi9sDZJ5hVIK6srCsUWn59QXce7
XlryfgKC5mWD4aUWG1/xjVaAAtC35VnqtVHdIa3HUb0Ne7FLetDtPuXoeye907D7
IgRq23D+yKNxQkEA3CZmJfYZ7lhLpCQmcZdG1HVr7NOZWnnY1nE3ZPPnRD8nfdZp
m7P2819/mgZYj03HMN40HcxViSbS4q5JSQLUT7dSQ4pwew3wdnsxoVraCaU1AC6I
5hWdgLH2ao3dzG7Ituyh53xUlE63eMMYjFEczsprw/CdATnYMsLlvXenzOLHRhj5
bhx7DnwbB7b3Mp+YSWoQb/4oHxSz4ChinFLp93fbzvldj8c/WQKy+2l2xHekAey1
/zGczib0FHJSESpoxhS/j6Ygpcav4F2KcMg1zmpicrVIUQJk7WLdK+DR4ooFnSzO
JYV732xoQ5XuRwNVufT3Pobj5iBRsQVtU/cbuUNlnNDyygKF0/082dMa71tkvEbi
22Fu+p1d9ReGAH3beiypKbKHYpq1mVRShFxpUyuNOtchwBo7UmvlZ/w9u+qSBWK5
lFBE5G7vObfnaW7xJGJoQQL+4NQ9IPoq842uFMN41tjgWGY+no8500C1fItcuxp/
b5Y9zZB5yZnz7HBZIAkc64WmjIUqZ4CiwBdrhAKA7fVR8Z4O/X7uDGt9S75U630Y
RtZ5BsuJU7FtJc1NedbhIJFGSJugb4/stJ8AR6Da+Dfegv82INStKTVPn1aFpW43
dB8E3vK+xHHgnIpnZHlKOBxZkqHvaP/A0x70Duass/XO6wschgOB1KoOXEqgRCky
6qXm/B7/p6XkGtWqK3eeLg79RrDyVIzwB3+XvxsCToMSIbwZCKYf/7YW9u0YAVqT
HCKF6fbOGofJ+MKFKIp+6Dy1BVXtS0dLub7oBo7nvksLnHumj+kzBGD1o3RQ9sQ0
bDqMgRAtxb99p2GENdS42JK+FoMD8fKN6JHAeBKHC0aRJnFiVmbY2SqKa/7wdTQm
7h2tQF5FFYaGEinpsm25HJoD+m67ISZ7ATDFA7DPZSJzEGE/ueTNiRpJVfn8VOV0
XoE1UD3JLc6c8cVYiOkbEyYTo07tuJ7702aRlS4cTh1rWmVZVTvJjKvnMy0Cb+fF
Rpm9npbd0EtaX3sfp+gEudtQhU/wvrd0/Ph1f03ZgejYvjFDcq3sYPslttacOSls
mNYxeng0YnpmfUOW9htTwu6Ul+fX7k/KwnxR3QyQMskdQ8rXwxfbx7kikHlDYA7Q
U/COB0IK9MtMymhtxCA4a5wLyj0zBIcwCaqQEScDRY2qICfo+u5erIc2lKw28EVx
/Yx9irM8luYQbZM0VBnWIOQ0gtsrasyL+dsRW/fDz+4HtRN3I4e403Df4wcrLzpn
FCt9lL7Rosp2Fwtbdo0Gt0gY61aRYdc0PemaeLsLRJ+kzKxGlqx6dkj9HbDaKh66
+GOEMWizbjtouRRA7yN/FcJukZPV1G7IpAeP2YZaP2+Atkb6334ZeexQ6kJqTQzC
pYYZ9XuQ6s32dpA0TwhV1rIkGEgZ+DcVL9JB/FiOD8Ui+286+CGAjzUulQLyoBos
aLG0/vwiH2GJ2L4sqKoBRfF/AIlx6z4C/YF0CqhdsShGPN1MskGCzM1Vv/S/xPqi
wUVWfHpNENsHFEkAUu9UyWf99TEQBP8b9QmB4Gko1kZJjvohaj5YYyAx6hXPdtsK
8S/QGpAy0Xas5NU2umDfFEYvm5td7nrWh3uyuG3U5+n6Ax49ivids8yPkZp7oGKv
vPaXKZy6oOtQdIzG4tVgoKJAQxnv//MRppVXr5LdZKlau7aFPtHudO07S8c2yd7b
7LlZ7BZ9OJiQNRa/bHXP7hCX9m2VKkP0lSLzLvacb0uGQz2Yua1tO1FOQhNx+Rlc
eKg2nRiJHyvGe51r0ANCha07URDefJ7RamYn+Ct/hXTJHdmAiSTTAmBOoPHfOvMx
svQe35st31ZV7XxcZWEyX3jxKhBe0q8Yn4aqs+uSFVcsPwArTY/VoiIbY8WJmDxR
sB75x3d+VDCJmGXFDuDnPKLl8RwRaB6tP8eqpY7DN6KrEL+Ngt63K74e3iCmTkxT
oFGMBr1FsqirJE2s3ss547m8z5honMLCDqdx1nAUKY8Kb6Oox6sQ+ZfgT7nSOElo
oY3C0CQtXWphbGYhqlf6NP/MM1eDJcYymxElUFzSZ7Ny0Mkw7LYax+QBSpzHz6Pc
4HZw4muQexESjYRBu17L2CYNUav+KeEXVkarUs/L5bpSpJ96owGfk8oV8Bk2rhPx
H+KusSG77k+vaXjWgXtVk+0dPX5QbR7cAyrRPdfblatcr461ddceljrgWX9TTfMG
Q09tOhahM3uBRj42mOoov1EZ3NO9RUcaPIX53bWDlrtFLxUCd5UgBIllzDV309Kh
Abn0EbwfB0xB1bJ1QqyOE6Fq3icUmNqXMEM2xbgd47x6dn3Q6FJNrsYfOMIRU61h
rG5c7bWptxkDtpi1+k9+aUAW1KVxfJTwJFUOq3DEuSn82lg+fBY2M+be9dGJHEN7
rXwsPWo0Xz04xE1m1ju3a5/RklKb6GqM8WTzrfMP25z7jp9It9CREBff944OMl2D
538eYQ1r3Oh3PdUS++XH66F1XY6b7i4U/JZNGDh8ToSJmzUSp10SAN7W1dw49MPT
UHZU8tr0+ou0TCyh7vJkRIiTAuN85W8ALVD3EkQwqxU0djySU0gHOQCNLwp26x/Z
YQaFvVUxNqQwP5syS1u+FlP0L1yGCWAiAIfJRQ8grrsfWiA2kvSRoJA4dV6gFboT
PjO6purewSTaadtkTB41Hj6DTmYHuI3vbAabA0IfWQy5IVLZExdpkdTFRvkwAZa4
yWIVncjqAwlfvtcbzrUQv9E+R++POCeKjGkDMobc+rv90Jefph+YxbKHAyRhtxWT
7LyjKa1xEPHGYaxm9dnlhpzS6okTnEqrL5Cu0K2jtj7KqCBrJsY7sUKGHLgBwb+J
UPKDE9HewsgkMB/M79Cup1MfExMoW6S+0cZWT/TuJJvxtufI0QUdt0noRmUSz4Rt
Olaqj10JFIINSRotylTsKLZIcBR7vktdLwBK9V/detnPvnQiQh+pCaIqfY4UwSA0
So2ySBy5OrpTSoJ76KBu6CAbKqX5Oph3ejlv8w/roR4bu0eg2kphcU4wm7lmGt05
51laVOhq36rhf872+XdfQ1mr+QCkRAIUTqpM61+Q8AY8yApsCYdIGbR14W3xrviZ
T2Kf5LJvcA+x25HtxDEURq8AzoGbXx5j9528oMq+23Rt5arhzSFO0/jVB4n72/Wi
IEeX3ba0N37nrnY9aXqg2yFEXilXofKvAtIc6eeaftRvVN54TUJ2nlFZScyVQtoT
Nd8lzkE6Cx/y6m6QzvrIuf7SFGDW8mU2ZFlqz5tL/yo14gLRszHbScJZDJrgo2Ag
9YB4E09YKvLQ6TEZdFc1E/s/qg60IxcNqqwt/7bqhnJ/c4EYKjmDXdAL3Ng+6Gei
lDva3wZM+7S7I/tRyj/ds5p5kVZqR1qxmkAWqNnpD1eUilqNyWQZrHv5Pb1P8W8a
+RS2DwAKKfeP3yvKWYG/X/ghEyfDXhtuiSKTO8xcbrU7rruAujvSIlyTkZa5q9vk
4gfWwiMcqntqrJuGN0LhWyjaPi02RFM8+NWWxukGbVw+NAvmKhctrXLGJgDPZXsU
/4YpWsJiwfk24Cec8XzA5ZpLzwS7yIOl93WBoHYU1zPwfpyCIzuF6/lvPGxovdkG
lX2kwDc47oWV/EbMuvplYnfdrw1YsPBR6OEEPRWCz6MAHqLnPVesvlTEGvC9alDB
Gf27wrJ176iEzGWidg5/XPGWNqCNonOn2xBTcY0f9SRLfMfYnJ+ImchXb1bCn99m
dptyIvalbyyOdpILWfmey7lTGpWXXVqclicUhsQLKfyG9FOfWC7/0IGjKCALWR87
f6qK2ZCxEbu/mMiunMtqZQlI27968wbRJQBkpVb9Fle45RdwGx2R9hUgDi2uLf8p
IF2UhaPVg5tJhiCbad5JhQLc0qLqkQ9S5/exSy98uDiHWCgnTNc7o+dsPf1aY9SI
6kvDEffv4QILczbzJ7Gw+NptUUSqQ3YmVIWjTHhW9hlaugH18xI8xF3KWXSEpbOU
hOmrrtYmbE3gLQHP2ZJ+ZSBpXRkfnILoQstBn0s2jzu6dVIlcgMgTtNH+8Nd/70R
CxxQLmktyoWhJ0DsYB0mnNXs0mLtLgbEW1Nysk2jID5LLINsHuLkvxOPPdf1dC82
RivrT3xd/PHqaGIkASk4KhDdcMzLR3Qfti6ggAYTwx7ExaYHaL7XuqKLIMI9sMRO
+vmJEOFetzxG7gGb42MADpoT/PHCQ10DqS38JDby4VRo/+mY3OhZRUrpgqGFEQ03
CNNAtwdBN8vqcTeY0EExhnaGVdBVuvTr3ttN5Re4pF/2K433gV1/ivZRHilWRQXC
UpQrtfTQJFK9G+AmXSjrvQHhnpPj8480IEyZ741XDEDli00ZKqExVB6gvH/3uBAX
EMgkAUQTKRizuDM/ThZ9o+yY3lnrUaaOjMwTf0UL/V/PkjHdpY7XnoXDd+D8dGPj
Rj5iJuXN8hkBOn4m4SLOIurp3CWQN1+BsP2TEuLxs/WvJ1mY09JzPLoaltc/eLfM
MZa19n74hVN9Ca4Sp2Sn1h+7LEyeJwlQDpvkBPKhopUPjvotXRdkuVgoMpssqGt2
RpWz/jy3DLdHjC9H3m053eilbAp0HDQzo419s/6fEyBkl9lZcelKjeXQjRRxGwF+
H6YkzCo9SPkM/9HSS6708Ciw/QHttVgePXo5M0YcDJpR/p6N/0uwGyVYQqdRYHJV
2rrUWNHF/zdE6KWCfeKb2bmAUz7vZg/9yysMNzzMRwIwog8dF3M3nFe+P+N2a511
4P16z0Oo+ZryanAF1eCXenkCsb+8m758MzAjSS91EXc2JTyp8KiGMdNheIov/DYI
ke0vIDfV4mCr74cRkE9v+ScIATrA2hHDhhbCBX12CH1P3erotk3pSv/6uTE8+VWv
/vMla4SRgzqYdVCd/7EOyJ2vjS4/wqYXj+18EM4WjXQ/rznPu3AepzyA9IhTWRS+
QDLhnziqBrURGXTk3juLrd7gyOkUtajgkXs0+wst89z55oKhmS1vYEw5mbkVYPjs
o0Q+f3gIh9D77TUCFravRf/wI1YlCSGDaouE9+3/OuHwYegwYwYqlSPlH6MGAyru
ICIPFNGURe/AGtdd1E2YxsaLqpYS1O8gMwCc46mm0ldUtn0/W0EyHZHZT7ZHIqKd
iUeU9qd5QRHj9+zJ5kKH3U80Px7rKEceHDEQsdFvRkNRs5K3D7pQhR4gy8Vox9c4
IreUkC5YKhG7LLUcobYustLyAUMVQjWNKHXTzKq6A5RmWzd35QVJfg+/gbYwuup6
OObMKjq/6WBuYHFZajOmkCRIVwPCGxB7MLrlRMEnaYYJxohJ7U21Ri3fL1JcOmYI
E063ZtrLpWCqpu9+hDpeX9Y40VEJSjdmNPzO4UEvf163Ep2i9VIGKr4N9gLT2WW/
lVqJ101fBitCip38L+90G75VrVYhUjg+xrFN/QXCMJqFxuJYpM3M2o0WjfsRZ0f6
14ZS/ytNhCmGiQqCZpBniAY5wk92ybIxxy8mCMHc5ZxCbEFWGRJOjgSG3VHktL9X
U4TysJl4fA/xVupjYcnxdiKaV/tjUsLqLmUs/gn256m4A34aEc4S6RaF+UdsffwQ
2grysoHMcjWoZxF7ltbBulFndEMXIq5McMdot/hBIhw2hjU2qe93ErfSAaa/Za3U
UdkzruinEBMhoXixDdtqIMjMsdTWeOOxAsevk6eXuiBKK4cbQsQyzgrdoEi+4XZB
fL4DYn+g87yQ1tu7N5SMKkmc5S2DwXVLA1M/XFWPymHF0TFv8F71KBo5TyndVlkA
QnSb91Q8eKCxmYaOk56NcskrIW/nBQsDFYkcQnKuCKYehVSTUe7DPqqCZTL/qoSY
1qwzOd0i6mGffS1WelBkRX0vxkbg1J9fNfz3eD9+DUiH1zcXHxqcDhljG168W4DY
m2t8SY3L5dMWwwA5b9A57EvMMXRccA8PFt8b2RIJWWzePw1u6lR7ESXbUXqTOE2Y
T4dWf3QgIYOu2s/z7rssPffTUPYrNwYmIy+aZsH4eCH+LHQI1v0uEiBfUpBAmmHe
yv66qHBbPIklCwGVb4uKK/eWiMX9mFWcqNcxG7+GvV0PNcCK9EvImQVwRiXonXAA
TmkEjGtsljl8oDogEG8qWD71tZJthjd42QSqgLfjT+1/1e15m/sqE/FopS1cXXWl
e444dR/5/WPbsyFL+zrTLA5OT+wFBpa0WqPp1mNzYc7BVtHVPHFdiWfB7cP0epeA
OXSnFM0vawSdjKNijhhoY6kmbZ97bd50yPT9l7Db5TnA3sGnsiCAGMCuPzm8lcgc
mMcRBP+bzIer/isrRqMYTj6Pvi9UcdM4H4oekydOPoK3Tbo1YJNL8+XpFyzGPMQd
iesRfn7CbJObaLUj0+L1eLb5yewgNMplLI66wcYvjcd9A75VCEqDVmLk+8FSrg9y
CjXfAWmfb5KQYpDMgObiDtWqWebA82xPpmQXurs50Sk5MJ+QpuSnqdcZlIRhh8RY
Euoh09whDKnexFVUsOK+354KSC0hGAmaixAGNIPed1UHWBreXfRvo/IklPKaW6iJ
6xWK/Y9fsTaRfiy3JOCsBZ1qn2bFeLutJYKEA5QYR7hSfaDjyCcd4y07mfR0Cx8P
axYheY6rh9xhN6OAW0FQotq7QafXOVaBKZChSPiYEJ+mcMPtvZI6LnAZuwF7vTIU
NqAAV1LD5L3/uNCyaj9MnR8kOtLjQp41PEaxwy+UkiBfNh5Jsr/bOeLb8RcE8f6i
wQvisnp2LF3QICNmlwM9ilVGRQuKo2FeqRp2NhCuvvRnOfRTj4IIHymgisbbfPSL
J+5f4o2aZke6VqJmTU14oLYqshp9AakM3DeNh1EbkwnfgEWRMup6ows4ngrwHrIR
7iV1O+/I9tLI2denJDbNXSGBK8OVVZJ7d/7Vm7rk8O/hMvvleIDQzRKFbY41cOwA
2+PesBu4d74zj5w59xYXJqZIjjNwp4NrMa2G2cMTLSNDleVWYO+WkpBBdBFBOvb+
mNuuJGPfQAFvGZFxnlPzI8dUW0xvPTFytcUizdCzzt5YuQjthjKXiDkxZ7si9xFM
R+4BdkAUs91HQNP1WY0miEHusf2K8/ZLtbrcyHdwrhNN0pjeVuaZhnI2yQ9yPIGV
bHcaVAdTTVnaK6HU4pHvJN4v/Jtm/r3UzWLvdvhree2A+qucc1kDmcVGynxODZVG
lrDwAplV32oSCHYIypMJ+tHFr4aPF1Qfe6LbPGZ8Rsug5eIGBUpdQnPZNVlKMJ6r
K+x1hNtin8S++6DdfOHgqA1enBTC3XdCHivMMRSPolHn9TYSkvInWxukd8UNstMS
2HZC/83sgxMl6COFFhhBd3tGd9IwLcq89rWzAFRcTkGpi0YzQGc2xnnxcxL7t0Ck
kEpSyP3c81DLYOnzoy6NZ94Inhfpcicb3dKkE2Fl9hagqPJq5ITPYCjxttET3NlE
yG4oa0aGc1pRVrSgAGThdm3zAvEUN3nUl9rQhsLutVWEafLx7wqZkSUNF+MafxjN
J+aXxhp9y5H4jZQdLXm3Wm/I7N4V66Vtdgf1dbSi6GxM2LXofFBbtxMMfo/NiUlz
Zjvu9qy2NkOuU9XemI4wDmTSrLIA2aHHACSF7OXTskDf0og7vutgf78v1W7Z0nTx
o/cQwhBeunFuneep7juGEiB4hoo8cIS2rppgiA/cgIFZQuXnUklImtAUrMLDa3UK
KVQi09p/ye0OM1Vq1UG64DlrAWD7MPz/VCtgKlbey4fqnfx8B02jKHIuaKh2vHQm
jclFJY2IP1OQzrGFC2JUyNyPYe8ys1eswjf+aBumtDlBAbn1eeRTyhTWxT7Ewmqj
JbTS+GVPzbDrmNB3vEroKuSrw4iPZR/tPXEBBQKu0Ju3CS4IlhtLx+qs37S6E+LF
IwM6xSeh/8JeED8kPDqyFqV4KwwyWzhHDr89ggUJRcbYadcEJ7e1xYt7oiegMIeJ
TDsvWw6V0W0iF3z6pQxOqyBmj1J3WWm+v3AT/OlYZZDJUcTmNrDTUcLTSW0aCngM
1Gmb0pEviLKtSZfvKV0Ov3tAfNMq5+KU4/JzTS7zt32bJRSWyNkT23IX5T4rpdvx
iQfF8Au1Vdcol8+n7EROfh7P1rcTqxJVtcT22zQpT67DJHNwFLr0LOZwPeFNctlJ
MzcLtXXhoBehj3mji2eimlmrwDNFAcpe4EtgJFKsI0nA7RU0ddhO0d2+Em4b27xp
EbvT5dVe4zeY0WKfXz8V8poeYXFRi43+oBHWBeEax6Ofv0zdyWGY6g8l2zNlFvSX
0MCXtRYeLCsrkppOvepV4gSFr62VvVsbu7pUcX8I1Tm/W6yV3dgvg03vjDtgz9oq
up85kYbQA0OZWDSj3OfLcOXro7BBmMQ76UJDMtOa8L7J2pxnH986VRvlmmu8QiDt
2bX/lzU6Fd6SO5CjhKrmUOERlRgMCWXqvbE9Qi8Cvx+hGCesUs9YtZ+dbIns4wQ4
uVKSbgpbS2j+C02av5Wo7jqsUehEJB0fUmC/cPeP+1h3e5NLn6fSIDtAcnwFYfvQ
wb47kQ2d6yE1azh/b4hz2cnh72vTT2Nj8Qi4Yqq2Wa3of7EuJh21WNzm/QoB8Sfk
OwYtv95MwJEvseUICc11el6uIAoOdlOj21TvEqAyUhhydWeNtqrMEdqlddN3ez7Z
ApZ15jzzOGjk6DrxiB6gxyl6JiU6Kd0863WF5ZfVcPsns+lHalCjwwoeUKpWv8+N
JGxrVDR5ThSxDmvCzjrsVKqYr2lLb906uyTXVyXm3g6WrxiZZzA3QJunfb9SGcmm
LHyEjT07uCCE+TAaSwZENe34FSITpU4EOKtVvUqYHOWIpjSMa6aJZ9mQ4Fq368oW
LOafhHQmFrZsiZQ1gsFqQPd9eG3iwdIf8v5inbgzNIRlGRpRRaPpVt1Is0PElblT
laiI/mWe4u1viuEXP/wpM6sWGHsE/nWKI379fZi7/IyiuD6EFjvh/qLeVqD0v5gt
b/Oe6+w9q/Quy/pKTRnwVhYVHoeEtt1aq4LhMwzQfo5YS1uMBo63VAMsfEdulsSH
1FqGIDtOF2zlJShgoZzrgaoIAzT+LNINz2Bi9j6Su8ZWUFkN8LkWvDnZ2hj0uQWj
Ld+F0WPm8DRSNNZe58UbmtqkZKBjVPOu5Jyc4GKNk2XybUtPwjMAVgGZYGladBSa
pKDTslZ/pKU/eOHP7juz0ZkHHsrnVWZu1gPCjKbXsZLBurFowypKEbQNKcYieXVw
XGPG0h4zIdgjyvWyaeHXtmtFIyKfqDFUH3yceon122IK7udLn2cyH9jGgGGhy3On
gSNYDEZu0ARb+yMlEXgGcQkkNua6xKxN/+AjWTRT+gxI+devbAVycYlG0CaZGjRr
J/zcTsIsEraVbGxb+iomqchU78vUDz/++Yt5R64aRsstQSYR7HrBPyk62rLV+Iq7
Gs8Is66oyMPWuD1b73m0ZpjyhwSThTHD7iJyQLo0dCkyFvjZuAtK7B+Ylxi3bcAx
AYjokZl6n2h8g9hKfcp37PNcUD60j3YgJF5Jfd1BbOlDI2bMw7fVoE7vYI9OZGhd
Z01X2PDGAT+HDN6Uz3aDwndhKukfb5GL3YkRHWHkcs+I4CQs/TFiEyR96mrd+Mog
+07/tK9sCBxd/gHEGvc7SgwIVV1BHXPj9rzIscftP1uhCjOxCpfj8cq/XnvM+Pm2
aLaYv6HYU4+P9/c8I3umNflRp6Sjgilz3T6h7BYtqVZb88kze/GJC+TaDENzyxO1
TARO9zbr+YTHed6n6shGKkvfeVVJmcn+nPLEieTKJFMSOVfY3Phw1axwBbeJr5Di
nVqF4jYWYqocI3DF7OGZpFh9Q8idGihjr3FRpWVufVgsc6uvECnjhM0Dxl0zGGol
kFGWcN+jx0A5TWeO6aJ59lBOJ3J2U5B846dKswn5rVa01QIFzPyqxg4axAPATRdC
PA79D2aBL3yYw5jPf5t3hhiik5Q/DR+hCnaqkbYjQjhGcd3LhT1UtW/a2tmyZKI1
BV/N7OVypYA9DctYhfAi1xRxbjl54YUr4HVDfNhuhtMV23OB6Z6qKWUaDf+ntsPr
uusdJY5CU0nolUIpoO3tn2mi8oINRgW096VANlhz2D6wEf9P+I46l0QN2MQLl/89
0mdzm15orR0zFr4rUDoI5mvUSDilSmLNiB3yBv821t95zMzHo91lT+Abv+BetmVf
rkha0x2yjX2yFAKsXB/u2OgIIHzf/O76rB9IpqmcxdnzAJqfGzoVdJWJWrcHCElf
bKHkggDQ3CuX1rMwkcJNlU1htu1JJzBwSySDQvjxZWy3XIhLcRQBZWFHHM5ApLj6
a4GzjgG1NK2E/XWVSpZVr8XaAKMVxLBy+7aVKT/DTZSYmUxLVV9/IHwx6gyCcoka
eXgVAtIsEHB3wPF8D1XEVyGb/J3D9SFELnkgSz9soFAv74hQkfYAwNbifDfizQeY
kKmeCPG5rmgkcOJXNI/9aXNrceK1LfpU2hRG+Tsxx/b8V+Bg7UxtDVUlr54HA+0I
DDvuByie76c9e0wlIYmTt29MwKsS9UBOlBJ5z15oWjFMM9FAUx/xvkIH+uqaiB5V
DA8AwKDD6lGpLIOJ9ajc2dRTR09y/dFCQTfBcbnii1iUxvF4wktSr/3KVBRt1NJg
4rqqUMRYsdA6uSGsRIiuOZ1t2gmycgwVcH/6+VtXYTI7OIh64MoQ41QpiA01aRAY
ombM9YCjH7CICykK3EdC2xqD6A7JSjRi0DStQvCD284KCqE0pn5Ds94f2EkuuBZn
OvUo2j8Tgey//9lD+embsK4N1aV+2nBKFuWrajNcOf7AA1TeSlQF51RMnD2x1f/t
cyY8KU/bMTpTBVz2QToiVvuv5EIV2xcXI6u7MXAV5RzaRDB1BhV0WG/E4vTBO5dd
7g/Dpcr9MpmrZPnKaXwXWS9ocR4TAjLWgMGjEB64MTipKTSU6+W+oLGd1ydNAXUL
WtRp3Jseg1AtocHiCO5SjYh9SPJQotippROnRvkdSVjN4VF5BGWC8m5GI7OgnLyy
gvEDw3yktTjOXdbv094OPCR3a9GdklvFX9wN9+udxe2H7LKBr7Qwr4hgTE1Axyo1
vrP3qfq2Lz4eZxkdqkKZc1vAUBY9yQgLil5ieOyWQD6VcZ1q3FjylbpIZsPMf7Aj
Kzs0+eQZ984r1sZiv4Bg/LY1cD+NUeNtsHJuliXWAg5K4Eg+nNJzfzAf/3wdBHtD
9BtjsnzvvsKQuQvwW27LK8fL0uxZj5+Xv6yQgh2QDk9liTti/qkgVQhyTn0WkWls
1Vwi/0hcVYJIaGXRRUd4Kv2PFyHFyi2LwIDY1vvdiGT1ssjiMJ+WHSbs50+i7L4K
mmph8XWdMTHNI6SgTdldz32aM3aZCGuO4uwvW2E4BuoEYhTm8om//H8vS6S5PUAF
1UYan9MqDF9l3PosN/+kZ5ObfPwCDCB7xTPpsMM8eoodi5mQKeQHgkD81a3BWKEA
02PUz53N3/Fv+2sR7EDGE45zLSo0dxd92FA+f9yUVc1ouRjKangdF3Vns9+R5ZIZ
mULsMOgWFbzqPOgwY0mmadlGozoS/dOTV+FzyIQvfhKf1kv3+sRmX1EoOvP9fZjH
b4ZXkA1JLN5QFINMuvwCsN2b60N76nN/UPQfjpRCtRhDHsI9RyUZXVUnpIzUc00y
zrfhm/K9V+HskKLLVIdNascpPxYodEZNjeZVdXTHOSgqkMbhHXSWxHFJ7xGZcf3W
QhFJyF8cC/+71rA/ykJz9bvHALK+3Tmah8zZwG/ko+Dhq1/rtLNOTG6kH1pJNVD8
et1xPNsrVTwdpg0MWk7mQB5jedF7n8jDcHzOlptrPqmZEfues6gwkVHnvp21Mil1
BvsoaD+zlu1Cf8pGZTCP+ZbsMOZGGn8wLt/Ar74ls+IMxRAUg6sD67TfoTRuiBvw
oNx/7YBeQoOue7NpsFEeIqiw8xGg8sIZDkd3XBHsF90816mPqWEAH6ut0IfqUQDZ
dhem/C5aURuf3sa0Z/o4Jh+CxTNXHlW0Bo034XBxSylApJq4kyJQIAd1oFUb1sPW
3Y39bUMigIu+a4jvZlv3rP34H4BozVkLO5JHDCNKi6Y462BZPsMwmH2XRl4aUVwI
inJe+jyrwMveG1RZ1Wz1H46p+8hiSqtEWe+NaQkS0t/EsBbxxesSOHC7/G3q89VA
FkFKCR4ynMyj1JK946uu27dS8Ry4v/U3YzzSaVeeFvyyzGUR2mdYZPvXuKgS5R33
1ihQi8CjcS+UXvBau9fVvuGUheoYA7xk+H3S8rk3gaGOnPTxJ3iJZy/HaNhamMa5
u5bv1TghIcALcks7s8bG8YUWWNkeq5gvh18WW2O82hy6SzR7jCfrwN1B8fKWtuJ9
cfYEBCY/Lc+Wf34K+hO/2DHRO+cT/GABIbjqo1KrcLi9E6JFRz6eHbcngiP3lwa7
KA9WpjHEA0MkDjVIg4nc4J2cU0oCCCPvUMc+Kca1mFGOhTzY4wSbq97QpUyvb7MT
QoGHlAWDxRMdsecGY/l+5+8X8CZXeOvNOm70xP9QKPIIXiXngaGp3hmks0WClIFE
DqCC4HcDeEPC19VhWlXy3BoPZ/LunmisWNrY3F6N/rijId+9DHLKYoZUEJPG4Aiv
5mcccRgTv83L2RtdlzERFpnJTgUAQTkMoX+QJ+JEgLNw9lY4KOuMONZSl8UOSYLY
wjPpUFOWlOohUxUiandTTGc4gEuhFT4hfZmre6OVfJEsQ/vzf5qRCbR7EZpqICf/
g+2EhpTUfaBgCknTDBXyl/5bkiHyeWJVBEWAIg7St7GbnT9UG32SiayWkOJEIAWV
VqrNvbePUMaBXeGVT2sSliBwnTWn4bPKemnz14cYVNzud5a0s/1nhRuf13+ZHe57
MSC9w+3MuMU0S2IXboWbLAaX/DjqPvJS1qRLg2lA7x6V3enx9qunZqc+cgLmWJv0
uIgAPqFmxU8TsBcoLBqOxx5u6vOsj2+ZzIOVCGeW6fo7FhxrCiuta94vD0q1fGBZ
qYQRKdNFlISALs/IQRX4NFyl503id5Fs3OekpnEm6fgoCbhDejvxSGEbtnUigplL
C9g2IWlulU6vpXhNssm1e4llwZ/eAHvHj7NNyekOI/ddSd7HkBo8Q9cw8GFlPS48
kCNwESAjVRrRV4Htsq5XRx5TZdtEDy7uqLY0pzvJs3qGjWrY9v6MXZy4O9Rx3Vf8
N/By/j4UUHfKJ/QybTfoj0wY6pqfjmg2Dj1dDY86Yp2iIluTxA9AcTePP5G5+iKP
aY+XrNrAE26XtyK4iOu+fji3oKDrOm4Op4c6ol14TEkycGF69BvSBrWns11mZTWl
LrIGJMtwxZWU3l+J9sTuCyk+a3gD7SsnzO7PnubYCClpSP5dcmWT07fB+ndaAaIo
lRCGq2shmLtxV0m2vZMG0AESqHLhi2FjuMcZe9rmVZhJ6G/nsWSmdXyFwxR4IbkO
19loGhMWAu9eT1xe17BHX/LXwZs0FSR7djpn4tHPiuUUNJNzjRwLC/RwoBCCWrtj
fHfhQgz//CaJbqedNZrXvq+drL7R/+tpVD1AopcfbWMJY2G5fsY4x7OFsJ7iJcPg
RDWrqJVDe0uKqpfDvy4YrXKa6CwNWqV8u/u7lH7CDxBOffLDjUB7s1R5d/mzpbZN
J3Aue03cLslBwm88Y1pUvk/xj4QNujfuQ1Vae+yB8vA7Ls+Of8xF7XKNwAFoLjIr
YQ48NrNkoK+J4xF432I8K/ItEGuj3wKnKZUTIVW0HUtNDCfJjkSW+1kKr2AcOZrE
cAH0y8JUdSYr6ZvvBaLJV99zGPbWQFJZ0/j8O3MssFW/f8Gnuq8xxLfQhO+uJkfj
WAEf3BYTREINs9vFcUzGZWPMwO7wG/TdjIkEmWcq4MiDUIox3g1C2VxIQTh6i6dr
SxDc7WMp4h6DzCXrZe/R9Y4mkc3oSwMfTFC8b1OXHoAwWlJwyBisRi2leO6RY+i2
qNDff6recBsYpczgNyUMvzIr/368G87fLvoP6KZrsr/eatq8YjvvfpckMfZ7m/w2
hINqcBov3C1YvFGO9cn1PZ7YB1ArkmJblJFzP4PfBcZ5assdD+zpTKe8eyAXZ8xP
RALsfrR5KFUl31g1bt5GCKIvpKdyo9ZlV53z5t5MW0gIDVNh/p9CC1ZKK0OhckYL
rOESYljLThK96vS4jGvUccEYoJ00tSMcW84gUHM/Con7J/kKncDWVXAPOL0AGaPh
P6jUtTbsukyS/ZraP8hSPMp3xRXdugxB/umcO/7x2NbWYb0fkt4f0ABwoK7Ddv+2
oCLOSDpf5jw3Imxi5AuD0T0XFdaum8STDIsqU3KSRSBzCu0RQAas/n3BikskL/ec
IdyZR4bxAYT35OM0poSJl6EKGZydpo4IT+5PNN+5YokodsAIrCv5FjCuw9t00bgI
8FRrAoD5aXxw3rfghmr7KrUXxFQUdcj1fePb465Tmink9XrPYK1wtc+TC+RORG2O
+eGP1JYnOL1E+n4iP5vcH9EsalvTZh4FO6RHyyh6oAWIlLY6SEvUz6StP77OmLDf
2uD0txnZRb2ArElm9P1MdwgkJf+KL/nS1Lfu32Gf8izm2XYpT7OYWBNMZ1DDjM1q
XXnx3a7Ryj6SK9QP1bsPc59LvnkUhz3Y3pcz8CQ2cj3ezrycWeWFQ45sK2OlfEc7
T6oRSyvB1Vkfk8Pa74wM8/nM3FQq+dYulCkj+w+Gnz1UTZNWl4aa2Ua764jP60q3
yya4NCL7GT2Q6uerYAmdxIZT1+83U5NhmLKLTPbwTFH3SzQwtIyULs9Ef8wgf0xg
ngIm2J7X36pkU32tIe4sXgUezwR2OiXKmV+vqGIiUbTx+g5G1tR6zcB1tJW0Lyny
3oC7N5jIKd8+40xG75bFo6cj/9lDcxTuWr1ToxXlfc4BXv/Ja2LAG+KKKCvlnWQa
BqRLk9/33lD82VlXOtLnPuubiWrmwJ1drirJQsWqiELSG89ux52MQlRBVAkMrrEw
JBqn4sPPkrOVydW3wxuK7vYHfy7w6gPXPGwnk518KuT9Kr2SgcnLW6ADKdUKqGNv
sV/So/PqgxrOrKTGDpYYKxiMkc2OV5RbOqj7LffoyKrOLyev4OICDHZXwcCpJr1w
MKmP619x48thZWPkB/hYKQpCiVTkdUVa/+mArIFW1zrYZGjNiGQDw6WLh9XW+yAf
fikw2DAcxJ3ETq5PvB2XlJRwNBcHSGbP9U+eEmyx8H4/k9fC70irqHPrEsNxQqSu
dNQ4nuhideEnEEIgk/bda8/rcxa6ZAgFoTIYBjFVPMmR9Otf+qcyXmdzOcfb5+md
M3VnkSSdX2XBFmj/XFKNlQ/fdjKbbngmfAKOLW90caAWCc7BFUTWyDgj/QXTiPRR
8khFD1wcfriwlpbLJiFIhiXZ6dcrovCsv5kptZVWO04W49DtRaFlbP1JlE+2GISC
C1nvG1n/AJyUtVtc/8dGaSfPVEv+98fSyfztX5EwYw/HyiGKkdf/LMJlzaO/lG/V
x8zg0twJegYYmA3uoEBEuhrgwkQiQv4JiYds0bJ19h7U5sFE+Rmrv6lfan3M4SVB
rd2WogVjfWIZKRv5pBFmG5/roYa20MJzPUOk0da2St+gfKYdDj7iVIlpNYATxf8I
URk6xQlGs7BPUZXFpo0Q33awJCqf3cd+H54oIqp0TT26/DKbvuuLinLxhWVAt8yd
MCNoBBXb9lz8U54bqP6cLRRvrJi5XncLWioCgY21Maqo2xEC7NWszmwEUtnetXEy
eZCThlFUwoVVh1sxn3lybIQnLasb///Vo4kwRpn3JVA=
`pragma protect end_protected
