-- wasca.vhd

-- Generated using ACDS version 14.1 186 at 2015.05.28.08:37:08

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity wasca_toplevel is
	port (
		clk_clk                                     : in    std_logic                     := '0';             --                            clk.clk
		external_sdram_controller_wire_addr         : out   std_logic_vector(12 downto 0);                    -- external_sdram_controller_wire.addr
		external_sdram_controller_wire_ba           : out   std_logic_vector(1 downto 0);                                        --                               .ba
		external_sdram_controller_wire_cas_n        : out   std_logic;                                        --                               .cas_n
		external_sdram_controller_wire_cke          : out   std_logic;                                        --                               .cke
		external_sdram_controller_wire_cs_n         : out   std_logic;                                        --                               .cs_n
		external_sdram_controller_wire_dq           : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .dq
		external_sdram_controller_wire_dqm          : out   std_logic_vector(1 downto 0);                     --                               .dqm
		external_sdram_controller_wire_ras_n        : out   std_logic;                                        --                               .ras_n
		external_sdram_controller_wire_we_n         : out   std_logic;                                        --                               .we_n
		external_sdram_controller_wire_clk          : out   std_logic;                                        --                               .clk
		reset_reset_n                               : in    std_logic                     := '0';             --                          reset.reset_n
		sega_saturn_abus_slave_0_abus_address       : in    std_logic_vector(25 downto 16) := (others => '0'); --  sega_saturn_abus_slave_0_abus.address
		sega_saturn_abus_slave_0_abus_addressdata   : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .data
		sega_saturn_abus_slave_0_abus_chipselect    : in    std_logic_vector(2 downto 0)  := (others => '0'); --                               .chipselect
		sega_saturn_abus_slave_0_abus_read          : in    std_logic                     := '0';             --                               .read
		sega_saturn_abus_slave_0_abus_write         : in    std_logic_vector(1 downto 0)  := (others => '0'); --                               .write
		sega_saturn_abus_slave_0_abus_waitrequest   : out   std_logic;                                        --                               .waitrequest
		sega_saturn_abus_slave_0_abus_interrupt     : out    std_logic                     := '0';              --                               .interrupt
		sega_saturn_abus_slave_0_abus_disableout   : out   std_logic                     := '0';              --                               .muxing
		sega_saturn_abus_slave_0_abus_muxing	     : out   std_logic_vector(1	 downto 0)  := (others => '0'); --                               .muxing
		sega_saturn_abus_slave_0_abus_direction	  : out   std_logic                     := '0';              --                               .direction
		spi_sd_card_MISO                                           : in    std_logic                     := '0';             -- MISO
		spi_sd_card_MOSI                                           : out   std_logic;                                        -- MOSI
		spi_sd_card_SCLK                                           : out   std_logic;                                        -- SCLK
		spi_sd_card_SS_n                                           : out   std_logic;                                        -- SS_n
		audio_out_BCLK                              : in    std_logic                     := '0';             -- BCLK
		audio_out_DACDAT                            : out   std_logic;                                        -- DACDAT
		audio_out_DACLRCK                           : in    std_logic                     := '0';              -- DACLRCK
		audio_SSEL                           		  : out    std_logic                     := '0'
	);
end entity wasca_toplevel;

architecture rtl of wasca_toplevel is


	component wasca is
		port (
			altpll_0_areset_conduit_export              : in    std_logic                     := '0';             --        altpll_0_areset_conduit.export
			altpll_0_locked_conduit_export              : out   std_logic;                                        --        altpll_0_locked_conduit.export
			altpll_0_phasedone_conduit_export           : out   std_logic;                                        --     altpll_0_phasedone_conduit.export
			clk_clk                                     : in    std_logic                     := '0';             --                            clk.clk
			clock_116_mhz_clk                           : out   std_logic ;                                        -- cl
			external_sdram_controller_wire_addr         : out   std_logic_vector(12 downto 0);                    -- external_sdram_controller_wire.addr
			external_sdram_controller_wire_ba           : out   std_logic_vector(1 downto 0);                                        --                               .ba
			external_sdram_controller_wire_cas_n        : out   std_logic;                                        --                               .cas_n
			external_sdram_controller_wire_cke          : out   std_logic;                                        --                               .cke
			external_sdram_controller_wire_cs_n         : out   std_logic;                                        --                               .cs_n
			external_sdram_controller_wire_dq           : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .dq
			external_sdram_controller_wire_dqm          : out   std_logic_vector(1 downto 0);                     --                               .dqm
			external_sdram_controller_wire_ras_n        : out   std_logic;                                        --                               .ras_n
			external_sdram_controller_wire_we_n         : out   std_logic;                                        --                               .we_n
			sega_saturn_abus_slave_0_abus_address       : in    std_logic_vector(9 downto 0) := (others => '0'); --  sega_saturn_abus_slave_0_abus.address
			sega_saturn_abus_slave_0_abus_chipselect    : in    std_logic_vector(2 downto 0)  := (others => '0'); --                               .chipselect
			sega_saturn_abus_slave_0_abus_read          : in    std_logic                     := '0';             --                               .read
			sega_saturn_abus_slave_0_abus_write         : in    std_logic_vector(1 downto 0)  := (others => '0'); --                               .write
			sega_saturn_abus_slave_0_abus_waitrequest   : out   std_logic;                                        --                               .waitrequest
			sega_saturn_abus_slave_0_abus_interrupt     : out    std_logic                     := '0';             --                               .interrupt
			sega_saturn_abus_slave_0_abus_addressdata   : inout    std_logic_vector(15 downto 0) := (others => '0');  --                               .writedata
			sega_saturn_abus_slave_0_abus_direction     : out    std_logic := '0';
			sega_saturn_abus_slave_0_abus_muxing        : out    std_logic_vector(1 downto 0) := (others => '0'); 
		   sega_saturn_abus_slave_0_abus_disableout   : out   std_logic                     := '0' ;             --                               .muxing
			sega_saturn_abus_slave_0_conduit_saturn_reset_saturn_reset  : in    std_logic                     := '0';              -- saturn_reset
			spi_sd_card_MISO                                           : in    std_logic                     := '0';             -- MISO
			spi_sd_card_MOSI                                           : out   std_logic;                                        -- MOSI
			spi_sd_card_SCLK                                           : out   std_logic;                                        -- SCLK
			spi_sd_card_SS_n                                           : out   std_logic;                                        -- SS_n
			audio_out_BCLK                                             : in    std_logic                     := '0';             -- BCLK
			audio_out_DACDAT                                           : out   std_logic;                                        -- DACDAT
			audio_out_DACLRCK                                          : in    std_logic                     := '0'              -- DACLRCK
		);
	end component;


	--signal altpll_0_areset_conduit_export : std_logic := '0';
	signal altpll_0_locked_conduit_export : std_logic := '0';
	--signal altpll_0_phasedone_conduit_export : std_logic := '0';
	
	--signal sega_saturn_abus_slave_0_abus_address_demuxed : std_logic_vector(25 downto 0) := (others => '0');
	--signal sega_saturn_abus_slave_0_abus_data_demuxed : std_logic_vector(15 downto 0) := (others => '0');
		
	signal clock_116_mhz : std_logic := '0';
	
	begin
	
	--sega_saturn_abus_slave_0_abus_muxing (0) <= not sega_saturn_abus_slave_0_abus_muxing(1);
	
	external_sdram_controller_wire_clk <= clock_116_mhz;
	
	my_little_wasca : component wasca
		port map (
			clk_clk => clk_clk,
			clock_116_mhz_clk => clock_116_mhz,
			external_sdram_controller_wire_addr => external_sdram_controller_wire_addr,
			external_sdram_controller_wire_ba => external_sdram_controller_wire_ba,
			external_sdram_controller_wire_cas_n => external_sdram_controller_wire_cas_n,
			external_sdram_controller_wire_cke => external_sdram_controller_wire_cke,
			external_sdram_controller_wire_cs_n => external_sdram_controller_wire_cs_n,
			external_sdram_controller_wire_dq => external_sdram_controller_wire_dq,
			external_sdram_controller_wire_dqm => external_sdram_controller_wire_dqm,
			external_sdram_controller_wire_ras_n => external_sdram_controller_wire_ras_n,
			external_sdram_controller_wire_we_n => external_sdram_controller_wire_we_n,
			sega_saturn_abus_slave_0_abus_address => sega_saturn_abus_slave_0_abus_address,
			sega_saturn_abus_slave_0_abus_chipselect => "1"&sega_saturn_abus_slave_0_abus_chipselect(1 downto 0),--work only with CS1 and CS0 for now
			sega_saturn_abus_slave_0_abus_read => sega_saturn_abus_slave_0_abus_read,
			sega_saturn_abus_slave_0_abus_write => sega_saturn_abus_slave_0_abus_write,
			sega_saturn_abus_slave_0_abus_waitrequest => sega_saturn_abus_slave_0_abus_waitrequest,
			sega_saturn_abus_slave_0_abus_interrupt => sega_saturn_abus_slave_0_abus_interrupt,
			sega_saturn_abus_slave_0_abus_addressdata => sega_saturn_abus_slave_0_abus_addressdata,
			sega_saturn_abus_slave_0_abus_direction => sega_saturn_abus_slave_0_abus_direction,
			sega_saturn_abus_slave_0_abus_muxing => sega_saturn_abus_slave_0_abus_muxing,
			sega_saturn_abus_slave_0_abus_disableout => sega_saturn_abus_slave_0_abus_disableout,
			sega_saturn_abus_slave_0_conduit_saturn_reset_saturn_reset => reset_reset_n,
			spi_sd_card_MISO => spi_sd_card_MISO,
			spi_sd_card_MOSI => spi_sd_card_MOSI,
			spi_sd_card_SCLK => spi_sd_card_SCLK,
			spi_sd_card_SS_n => spi_sd_card_SS_n,
			altpll_0_areset_conduit_export => open,
			altpll_0_locked_conduit_export => altpll_0_locked_conduit_export,
			altpll_0_phasedone_conduit_export => open,
			audio_out_BCLK => audio_out_BCLK,
			audio_out_DACDAT => audio_out_DACDAT,
			audio_out_DACLRCK => audio_out_DACLRCK
		);
		
		audio_SSEL <= '0';
		--sega_saturn_abus_slave_0_abus_waitrequest <= '1';
		--sega_saturn_abus_slave_0_abus_direction <= '0';
		--sega_saturn_abus_slave_0_abus_muxing <= "01";

end architecture rtl; -- of wasca_toplevel
