// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F5YDV3eN+7qvgBH3+fv1PuPOKCS3q+6CcUoHkAZlL+ZlbcQ/Wy2fkwy5s4P2DL0i
C0jhBpSLm+2FGRUm3DqEX6mwXPkBwW3lL+tN8WGpkG+DIoNXL6L1TM3CU+z0uaa+
ufycjig/PvNmGG5ZAyFMtlqGR1S757cIcHR2WsPDC/Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
lrvQvjQlUOdQtPvhb1aLlyHTdQqb97qquGd3XgpI9+j32dtPKeBxD6E9rBihNY6o
BFeQquIN9rm4BJBQ6sZ8qYuW7sfUVBrI6Vq8whN9sQjAjvRfXzbwf6T9rWckBMkh
L66AcbCj/SxgjYQ845yx1r7MFQyo2c66y+XLkLKGj10nZDCJzRi12AqM+SRKKiq8
phnJKYvR6QuoYSMz4K38+JLe0q79U7ntvXHgM2FAoQ+2/PcEhjpJ/IRv2ghEGQoU
ihrlsbjXVy2BrCVvLcqy3kLgxB4YigZZkBjP9pkaixqxd3xXwlMwpC7R5vlWquSx
jYvu0jG3wAEAudzZC4/VTRN4NuHU2KDFTqE3h3n8dgq+W3Spk4at+gdSboeiOimE
x2yjpidi/KSUe3vshW+pFieT5c3fpdr+V36eHtCeZ0FzfE/1pfw2TS0C6JzdcYJS
C3comC1rGJR8OZgo6856O3qQyZ4LRmXdmgFQQ3htvIJQ70zFY/WLin8SOYIdZ+Z9
auMNsBnFUQHf3OIk6Ejzp2HmKVDdBDVHhdOcCq7B6uuCuYVD+xvAC6SgmWc29m3d
BjJu84QWo19S7+Y679n4t9TkLjegmzm+yO0ioxc94jlcWHAqX0y8LJfDi9TuYOrc
ydh5FsK/8V7yOwMtE0c8qP2bRiFrmzOEcb9LUjfKGFuaVjIgzgi0SSpwZ8RwYD4P
U5K4VbHz8rpC2tyOLeCsZd5NFatzg6CmZ20UouHxyBQWEl9Ig0XBZv8MZ+2tkmSJ
CL9L2HlUB1/x41yJRtn/TqfOC3FYKbldG5OPIBmrQ8jeOEvhwS83XaMUqAXM/kGY
jKWsOzpXnQU9fyWGnpLZWyx9d2wKMI0JoD6jJhX0xcdbKGTyhA34PedlRJhQz54a
6vC4TVx2rSeuYWamVkryO7WLqe0gxidoJVsMHA8dLLFNOVNK5fGzaD1P1x4Ndbtu
FDd2BTkbiEHpYxHwCga4+8ogdmL705VPWiLylRgCGM2Z8BHhOzIJ8vCjZeR+hdZf
O1F86kYBQXpvDsfs7zOuE+0IbHVfOCKdCTBtpG6BGvl4G3OEAMtQbKV6U5JA0HRV
QqlvNYSC941HZAyhSKrJOqW2EMfvE01zM8YdgtLNvP5IjF4ZChBd7sqvHn5ICRJD
+GsB8mtLcvip5aAVYB2/+IXZIk4Jyeqnvsw9b+qse6/oRAC67NYDp/0u/TK01XhE
PLBFHboBuK/0nDAa2mLIPffj36Eq0pwsJy7vv2icvcUZFFfMYafaxTsADMzxsQYd
eRRJ5oDrb2fhbT+Lnnmoi7BfyDJ/QXQVgt6cI51jWLHDHY+sOmBVjzz1pdQbouG2
z5p91Jy6E/5tuSaJ7vapxWmEvBQa5D5gwH5JUgEKlQHvJPxLkB/n/5+5H02B3LHS
ChzpMdN2RZsiG0vCrWZEUg4foc3Ym/QhJEt6wLO6C6aDIHNaqXGJiEM0vs7jPQq+
NUD6hN39UYuyglqwlivKEPmYfFCfoj8pj8FcAXbmwtCQuD9M/wyEiMNnca4IIhgx
f6FISk/0MBKUv/9XSlpD1cQFNM6AZQXWPygLI5oh6bXhccwrerLcucCbWib6FWGV
pYLOgsbuvZ5DS2Ci2FU5Ku5ihl0uK4YWVc6uEZu7sP3xHrQ3XI6LX3BcVP+dQM/Q
IyDNaQutjWnCGRUgUIbNX7XW5X3WP1322gAcOaRhgTIYMiKNG+perMLwt36Xf0Jj
4ZWy7mN5TuBeOK4OcsKz/Iz7odbTEF+f/DKB6DHZr9w9bcLYpA8fwgtiNMIERtnd
LDVhD6UEsVlTrH+lbpfwhs9NcO1FxhMDI8NHDW/98UNhUdnw4ET8UAJwbIucilZR
1DnHTLrcdZLKtqWu7lYkobLyhagctd80ZQZqQdVyc42YBhLHH9G7JhKz4OMASRkM
5VmkE9ZNV4SvP53MjldFN8oVqD9ynxDZzzmjhfRkWzGi5bAjm+TFK+j8bE8pr8ne
SgOJTAlCCK7Anwe8x0wDnnGWiSlsB7hTf+E9Kmlj/YHxwwrvjuQ5fQHVIuZAnPlQ
aSFrYK497Q600YYOUXfooXsKBwNYRiHAZUB2LnGq+myOMcGMywBvkSYCahyQ5L5T
K3W438G3yXiztDU1B7f+/l5Ihso4tlp+pyXCSZiHAJoRQhIfhIBOePigOU3cFzHg
QzEl0m6784Ed+5DYRVk9q5Qn6fFD/OSv5z5zUMI7Y1UZEyN+fCVguyDdrGysjlS5
Yq01zI2DqpacVo832Ck3Y7JOM7hrtA6LyJNEdMYrAjBTGioyFMFoOjar0hT5NAX6
D4dHYe4usX8EZkt1pwsTUrNkx5+Z9s6yxeE07Q8yIAc5nTo5zuybQECkb+Rkqsw5
k7ZNC45MarLHg7m1Y4U1Lg/mkYQ3+iTwMw1fwDz/L7mcXIckwrP2+4m1ON/ywoee
ruUT7SAaXaBtUJTVrzVLEwn8/6IwJLW/CBZoPX/m05caashguHk8G9EU2gfxFUMm
uQJwlhAOxrndRategZy8zr8/XPdAd+MjIaRe39PMjcWLhqRthPgsTrTMfXWiK0/W
4ZzrAmgQgAhZh0SaFGWMokBie4ZM/lwCIsnvofGV5gp6PK/lMkDwSgvN1bAYkV/6
bbSwks9odpbDMZVgaRrH3wTAy0ssPD33M4NhAqvm5Hubaol/wkoaU5QjH57GAoe5
Ks+uXFQXLiwj8iZcT7S9X/0RWLa4WCA4ESqFZ91QyKFl0JZ1G9gC04GKscM/OLIr
a8BOkOJKHyMVnaVYv9x0xpAzYbztNexlGEAK7qxifh3exdR/BEKgTWD5/y7idh8X
MdVbOIOmb2Xm51milZC5uSJgr6K7+zo71q0HjwDtgnqV69db28kZcCFA+PE0zhvK
tGQo/4ZpmzrfhxXBR26VgFRVV5w6S602TxmRDmAivW/+sQ+8DAA1pN49EcXjhi3F
sE6ytFCITH2o7772G1130J/7fbdTmX2L4D8jDmPcTRymWhx8bjoMswM0exU3wIsG
bnVJUl4YbvM+JfrPNVz4+12qDNKE7GfhjZYDSnRHR93yAGX2QquG5O8/PZeY4Fa9
R/5pRUsq6oDIoDRFRWV4uiAi/Hk7gyVgvRPsb6VmuFj0Ft+UO/x5vu6gHEg/HF0Z
e4/XNTvP5vVoKGoLjHM38gBaQpDzcyWja87nh1F9SQhG3IIotDp2MR+0xzq4/42Y
+SeKjFPTHBfdZfelvRvrfFHbN1nImnO3iAvI9GHm3q3Sh9hKSB4wwoDYKGzhszEs
T+NSOaW8Go9XTdBrLvlqBrqt60ZbMZ7YWY3n1n9jYFXJRBKmq4P2QwHXUPdDhPzU
G+TZoMxwa2NcI1REGvY7SpdtWPk065PVM8FTRdVG+dkIOy/W8iatFLSKnLq55aiW
x6x0gn0c9TLvI5yJk64Kcr0bkigep9H7aOw/1omJX3coNEnPJFqJdGDVsiXAIlrl
MW/ECviqVaq18Iw7RtnSr3kc0TyZUcIPdliNNEw6NdQFmloM2clLG61s7I7Yww2z
e4StoAoN5/UQWw71u91q/jJUqWPxbLyeoNOanGicyOHSHGHRKu+NElwUNcUfFsXl
VnBcfCQvapyFU1ZnxPHqzE89I6OBk4GyWWYUOxbYSpPI+E7mEwKeSIATeXgQMTNU
iMZMjk9iSVIKkj1PAqDO4/pMGRDlP7/VMw8sXqZcscfZpBXSxx2EIR8+WB/u7kgY
jNIXK5gE99qtC5u96uVQCK+mNNr7Vt6WsPEgkTeG9gjF4Kl6Kgal8jWz1HDH/c9S
HMSS6O/UBIcSv/O3ntOZyt1+6Z1TdZE+TpbsUPO+1KlNVqlOSvgAAfYeCcwNbosL
AwE3OK0Mid9s88Ds8bHpXOx1C20iCGy+B64O8AWIlvFNyjpJPV8Uknyxl1lXf0rI
MmTsbkWeFHNNADLTg9bDosmi1yWjzTBzBhFiwkRM851XYlin0i0Zu/5qD5IUudtp
A2uWLr9eqzBBBKobW0it+O1cRRUSMAa3rkhMXqr4ohpa5HhCwBwS1cE7DQqx89kG
WH1bhS5NDZdNSfa3cAKQY8UYqQcvc3Th3O+EiSq5YI9DiUDqg3Y9UadQiY7oIPJs
qeHkEYvmt8xtCbcqKy23KiSlQQjDkn7uOmWAycB8oPo0gIyzns+TAMe86ZUzLf6P
4sMs62MV5ib3aBer3curv1DjLYr5Hyy2lRqwQWJS/SAwiXxS0v8y2CNsnb++YEwh
YxhYoAL5X3dy9bfIJTNqkaqj7cdOWOnHmiXrAVfKjn9yg2Zx8l3pn6KuveVTzyJe
w2HNJ0X62hdZx8wWmH9rde20GHdVu9j3oLyS791Le3801ff8ssfgKxsg/Msqs36W
43iLJ+qdPRqPfdRhcTZ6/cnxfdl0c8I+snd2Ea7XU5BXRxi6Qy6afsd4eQoeBsgS
9l6ZdUddvMgrsjN0MIOoV83iPFFOLIoxU2+A8AMPoOg4sym5iww2WcFyiUb+wRX1
6VKjj/tl4YhBBrDb7xLoqYGeuHHA79mKPsbzhuWWZrlJnke2hmeHskpcZri9Hh67
4kKaUNDLDTYXMsnuQieomLZ7SOJYj3ranHI7vKzYu4YP+SVTcOkPY/X+PQvt3TqZ
o+foWL+FA1SaGpfpt64n2GmJXmX2z9gR2AlwgNdlJsqaLcK2OGWjPgxhM6CmC0bG
UDy2hbwR+si68ZvaoELpeaWDXYzwBhzxq4PVDqBV9t3HCjc23VMH3XLbipJ/bRHE
Zfbd5NN5WRtMaBC+zmpo4cTxu/i8LaXQK3sMd4isyfsdRpAvNOSlADIsP/mv6/eS
97FABL/LG4g3Uc2X/b58qai6yCcQQhK2KbtVGhBvfxv/l7KxKQBTPOAfncI67w97
LhxbiriEDOYNcgCHRsANoDGjHnJh2T31XDWbol72+VzywY9/nUE1SNO1H1kN/pwL
UpJCsTHj6s0ujxc0HBcHL2OopVjNYgfUC1DXB257tYY5gZQF3uZGYRaIWO+0mGlE
4I+XHShDHAoeIHr7vUXbCBkXEGCSzKLlo/UtTdeCzOJhR/cgFlWy4ssYnU1ruKC0
+1RHAgwY7QJ596IWLpqoAVMbNoTsjhIn7GA3GdeEn90mD9oH8H96wJYS/xD8AyPg
AaUJrD0Jt70rdrFEFK+AlDIULaUmt9kraMepcifNACtlByixEk6qB+tEcCIJHxe8
h/aJa0HybRD0H7Rx49Y+AAGEshA9KBDj993ozXPf6cS7iegmUi3X02yXLRAhxv5D
/1vrEyureWCPOBzG4kSOiel2F+53FvmcKrqnVojHQsLTwJVf4WMlXiIuvXS62p8l
76j6iomp9CweVoCEGM8McaSHAOnnhIXJ4WQ1QHRBvfKnfbfu1mTyq9+Dl4CBCkSk
qFN2Yk2qhNmT3+vPHCOMtJxBsXkLoqMNTX6hC0XoaRuxIcZgIGCBNyqgyN+qr+l4
0hcong3x1ApeX/n97X3P6CW+DnuSVB9UrTXCznJI2+Gc/9fA5ih5yAhaKllILUry
DzX16HMtiWKpstfhzGjYIUUu1IuwkBX80E+Hie64pXuWoj/hL0c+wBYs8laXq03M
RMaGonFd/lXDhT9vq4+aFMONkGlMW7LoVlT5Eq/ix8Lo3fA0m2rakJmSI+LuNcFc
9zh7wFg0l7Vdj1cNcO7UXpPZG31Bdj67p+nARExyZmV38D8gQGhNbDJ4ez1+yMpA
K9ezFO5hAJrbr38fugSSSjjt5cuP+TTR8X0JxKufdr+BVS3SgofQ0VFsRTVk3MX1
zNHsE+7E+OqLLVXzDh0gnkk6xxWs7HCBZXUSo3sIQ7mKp4HYU+CYkcy3Xnu9XbN7
OYFiJ9vaeOWa7uiA4iM6jufOAjxdbUiKRlUza+ZZUQj7RoNvfeMR9CIi1jsSXpVe
pXeQiG5s6EUgwsQ7HHSmgqAT9gNSNx86/XFJCChILeBQ49oZlehH6vVTClXWaya3
VycyQNgv2YFvRtcqXzZncSVfUsMrvznEQdb0ChwLezzzUFfordZrudrtcI2RLA5l
VVzgGNmhcaXkdf1qIfXZMXcIRSApMw4wpQwcnPjLn3g5TyEFo11leUjBXdvWBtvT
pAIUiN4cW46EypvggvZIHki5PufggXWa8buvh6HFl1lJknereoovkpH9WDGWUM+k
/BLqTMBCfgga2KZ6eCeu23zmP4Weh+ibM7w5AghlVZD2869zAqVY9BRy2vtbiEbx
X6eZUpYXaQZVs5MuSWj/lYgESVKOLE++7z1wp/pMQ3eAj+cpWp/E/8z78ubwBPXb
sXi1MXMmu1XJgWxzBMod97DMecdytTyhC9+4RxOjRgSzJJwzN2NgkKNii+XnIMRE
LS9nUhumSEHo/p88GmMPVwWPq6gttI5gQHUBXr8FMhq05EmIrIJD84Alx1w3iYR+
W8Y3kkYj3KjRfcK7hgkOuEuWdC+OfKjPB4pgpiSVca7Mo6RkyaOhmxUhEUQS69oE
SJHx9zZSa8tZgHrptKXpwKQbb0I07crI6VEes3jiq74RtcI5a1AgOrwVWO5Wz4yL
j3Z5EnvSgtBJbtR5O9KFLORIPx+63CgpC5fjak0d4BVz1InP9T/nlu9Ul9IJBxOV
iPQjsqKAMQJDmyaTcL2y4oOTzMXPE4ufDEco7jhBylyXTNxdA8BNt2WtXO5BeSiZ
HP59qoFWkUflbEaZhEV9QzyLGzAOsSoeGAYz1jEpuu/9k+z9oJTng4fKgcgewnrn
oNuzTz8YMhxyZtPtGebOeofEyLK5KMKAvbT0bYqSId8x9KQOoz+RaqZR8w7fwinQ
qQspmpXMOS3JdJ6SwaN4zn3fnXLzFkUt4izQy2SHAtYtOBwtY+ZpBaiQ/IdIPD3H
ZdrbzODI9CV7kIDdUx3Sy+hAA0g/eGIFskMA6A1CQOf8nMr36kQ0T7Bs9SluQ2gM
lUlHQJfqvK57v6ojAtm8SXAYPLAvod1d89Of8ll00NRzkItBRlJ6YKc5X0QDXWE5
Xnz/fXOzfHSgcWFCOwAfUPMae+MyBBEhF7x3imsLqlV5DCK5a8fJZKlU+7e11tMg
3O41hmrDcGBsQZyEy5SZuUGSrxyHUAQPcag7P4NQh08J3Fv2kZzGiqKjLX3whUPY
981MRUBtLUw1G+Ki6V6WK5SbHpxlsc1ZO1r0RGWsxGie1bPFzoJbzlFhxDhokR0d
un2qowTN4vZS1ctlxOZilinLkZ058yghTHVjZM/el04fS/zik2URnxFK6fh6m0eQ
GrAVNZHf0ZQYHYS8kxUw/hb5lSnuyOrErpIkq4ScE+IBIIhi4bSGarL9GfxW3UNz
BklfDLr7TzgBZWcsq6dl6zxwFp3mQD+Je0QR/6nm00W6ofMJAGY/NOfEFO+wYog2
yXVWutUHiLxqjCeIveRRyhq2i+d7rB6xHzD+bZx67Wz8+AATReV6thjX+8cAUzo8
iZ+H1bZsB+z+auaRtjpaH92BCiHcEek4zI/To6LVKer18CjexXsCAxsAor3Ys4Fw
cTwvVw9rvnEC3hXeGQLvyl1uEewg5qyv54SZmq6AHrEieV2+WJFM5JmkOcy3stbl
xI3Fyc0wEWAA3rLcX4HdWoLVmHRLtCXhvSqPhTyTABYKrHJghYwHoWG4CMj2qvoR
WVetdJ7o0mWcuh2KkMxWVzFYnJPFHyWM3vjSu1kPmU5eIyBWerg2+8+D6nMmyLH9
RGhDK+FJkcaF0fQUEf2EpHQNRLSHvPHG1ik400V6Hx+IkC2gzy7cVqQ1yfmQ7adO
GuMUSOR8Gu2pDQs39X1h/+peB149CH2H988uAc6mmJ/ACqmy6Zg8mvgfxa9GHQ9y
eWmQN3c/8QoGtyTLGD0ZneFjqD6H2Ko7Nn9eDv5QLHmhGilsCAcLwZClKM3PG2P5
4FraxIrEyp9HonpmFb6LQok0/HPmCheeQ1OE9CZeC+p4EW9kLGAFJQD7Yq+bXwnU
dQzmQ3zEC7GC9zCJNVAHlgAvXFYcAPlHodV+DNxC3Bw801pqhATyemt1nAxHVVoT
l6wrXbtubZVEhm2ntQBwhEVP8KDLxH97Z/ASSBJ7UZzp1VQ8rTjGalWHZo6Cahlh
kr9xeX891LKg25nUw05ZY3GYGAsDRCycjjB7EeAqq98+KbygUGs/1pF+JpvBBzKk
PJvRvVo+79GaoGH4T0m6YuSMdmUvusbKc1dy0hIiVTVJNw5+Ry7oIZlMUYH62Nhj
qLFcQDRa77wJOpWyiJyGfCIYuFa1zLCG/WpKBpt1m1trvrv3MHGFL/tWVzfpxTmV
A+Bxuk0KCvwa6Uvr/30dpJ3/sgt3cghP3QR3TFBrFW67nyvVniGbaz1CF/bTfaPa
igbIbVkAR+1FB1tnQUccDj50YOhIdhMUnUNkhzvqivRegKq75k0Zh2Aa4w+yFa5k
mSOst0dPrESuU20cLChxC2cuaEWTamVBw5PD/8YEWvqQyUXiPVxAMuntn6RnmBX+
e+V7VvpOSXpsp+snkSMRq/lhYvDUz+ikGrkBjQzd+ETvvtC7YanCEJtx7AOiQFgW
X4Xl8B6HxriUduvLr4YF6ijz3A5BwYEQ2YctiHyPtPBXfBWK9RD7sh/dV9hI0MnY
PXRE6I+VnZMD86ir9WxRsdXtMC45lOEwfACug6glxAhEF1szUAMMDOXUDeblGZKU
p9dTrImfUjUZDT2fkYVnny5XgQh5ZBazCyCwQr8Ualkqj/TUu3cgFgVsGT5rsU5L
ezGDA/iEMXW7t1cQUwxqypFB/yJjo++b4admDfdqvCsfiTVzNqsOSyrP12jQipWL
l06/EMLmZ0+kDiCLMITn22/8Pj8pzXpZWYOPLV/orHw4LGhl9cP5wNpIyHhMVypv
1LXct1ejQf0aIUB+XKvlJLpUEBL1e6PeAzp4jpwRxMsFKmS1GV3G//xUBVywslUO
qxH/gXkvUaWFP61BMccKReXQmVMVKO2qk/MGZab2HC06fDFmdlKiu+r3bjNgHRX9
MRSRVDYt/g9raprzuDl/sCg4QBiurpkgqdg3xX3UDfgm2T9++dCVUdDwW2EAYn+l
mRj2G95PAV1CBD4CJW7+hNcg4bxzefFimc54PbM0b/pkbzIflJ+0p5nXZRx4rWMu
us89617Y/pffmWJVOJ736bhna52pg3tmvrqXLVLrvPHgc/tm7jS1xSlt3eECSbiP
8UXgjNOXc+q1aK1aEi0IRyne7hfnDWUBzisiomB351lihaDGQTu6B6wPmbfM/oqr
tdq36xKsIvzxZRr0VbdxHA3b0AwBevynqv4QiKPCZqbDdPCWwGwgYkf8+/8L2dzx
45T6L+2cTYX3KL+pGEcdPnr3AefcCCOgtv2Aal7TIWmxCcBdIeywhxYUaZySF1wR
wGzF9UzZPOQ51l+JZuZHt7bzWYAcgg4pFBZs3WTo5fs96kogJgvyITFlFC8KrPiY
GmiCpVVgKkqIKNuCS0naa3BtkA1FkZbxJg+2SfN8poxoU8P9Q1WjzdQCmaRI06lM
KchPs1VJ7rsClQm4rBu9N//72E8eSJUY66Mqd4xAiXq6gwcNA/shpzzcsXZep2sg
zzwxTpw2URcWiBwbkmCSaXNJubkSok4QCCd0KzRZS+/oydkpJJARzQ/jlsHvttDt
QVhlKtaCTGYfWsyQVUzJ6mPGNQVk4S8jjULiK4Wyv1yyCka7lHvZHlzrZxI8ojlc
eaqdMz1u7yg9u3E//nfzXnfYn+7V4mdiefwIsoTjYZVC9hLYXlhcDofJ43rxT3li
9fhKoBq6FrvV9+v1TZQy1a6ErNQYyNIYvy1PFlDiyMFL4uX+eGV+h6Pq2vsRjFEw
arOXTIBuWLd4CzpHsM8XI7XMWrU3uMc/haDgpVLMyqNgSlupWFfXH7Dx24GOWhRE
DRGt7CB6EerOc2s7f+EtB3QbFW/si6Q+lTAs72S3GcNp7DAsAQTnmQOh3IjGHW7x
s8NzK8Q1wc9+VMLKLfWS4t3HMlGowWswuh+Gz23+sIzMM1HtLc12AMP0F82FtOak
G033hXTYu/y7RWlAf2H/qN/xVAeH3tDNo9ZbERHlUpwuAHpPFUA3vOHgGZqAO2fu
8JjN+JnIPpFuH/7mGJFp/D3MyEOLEBbKDHYjb7zDxWdyJ4lTTZgObXm+SzfOImFM
1NsXF7k56kyAgQvSJ+vTjOqlL4PRmj72QgtHQeDpXuIY9uzCysjGXmer/zGPeqsf
Pq9Yew5f1820JvSJ3SR46AqmPSnog5Bvg4uvHcoc/ngu+Q0s5wvaravovpaxxQ//
PkRZMVEFCVsMkzkkrFIBMuJ1Pga7lU1WLRVDNdAvrrhfW84IzD2oN0dFCwln9ye3
tX5fbfuHMxgffHoB23CT8kLL50+B+YWEFX/BGJx+zFKS5/v0UNR6Mg+P7WyZOhnG
xRwqljdoQPrw4l/evgf71s553ineUS0W0aoEaetQiGVOiqziDxnucTcTStYZ21V1
qcmlPHAPFxywTWmipbtuNhL7fmVqB6tycUmtfEx+alFW1VyGh/R+5N+6DcXHtBkg
wt1zfGyk6ii9KGcjH/vc9EvX42hX+u+93I2fT0Eoe5qKjM3w76FqXlAQ4iR+xTTz
XRjpnheqlV/H+McGdtmFZd1HgtZWDJ77s5sWNyE2QAn95ozbyk7EMa/BPoYONrar
W1imx8TgH4RSypr/o+esNzHKUFnGc52Qd4o5DIAVB256dAZzY+8p1Lv+W0Veg+fd
zcvpvzUc6dtO20qlZy+8hy6JH5B5EAcVVb8v2f7ltyPVp6WNUgVaE3SYwm32CZLf
57vKcC6GfSW/gP2P2KODzFHt1qu/28glWJzYeVuPChTmKzCfNSr1NrRMjGSdjdiR
Q9Jn2NRM2JbXH+Yd0MzVmSBEm5xfRgSEMWMlbUr/aB8mMkVxpveCj9g9UnlNvDHb
a2Qp5NtnhN/uJplLCsDHDMmj+RZOWJIFCc4QgT0rXxzcWT/bo9OOWw0Q5MN99BB6
7BwtANnMFYZPUsiQUJFEfZzaq4dcyK4TDTJ9RmvuemPjv1PRCKFWQpE7sVfo7Ouh
UAR27rXvXAF74S96oBSMUdixZnJkzIzxuHGaoxA3UoO8X4arkWE+t6t3yt8orvbN
buCgi4FuYSZhuBjDsJzSY1MEBqUcLVGuQG784/E6Eqo0agHXpfQfavKIzDswD2F7
BUpCA6hLbjJx0y9z+QCt56W3YIc9fCUcDncxUYSieFQ0ayuLBF+y4CYshLFNp/DO
BiLg8GCpyHYAuaCTTFL3A8/CKcw/GErTyyxafNeqz8lhw7JEUWxxRepCy51Rcrv1
SzVPvFBl558o+0/eGqIE+RPTTfx4yKeqaDZEjLrDcRLf7mfAXPqZ3NVCwtPB1U7M
bWACyx5GdW5vPyUQXM+s5kKqZXINzgzjXCemd/J8AUMS+KwTudNClz8XftzG1r3n
APP6b2yMv3Y8k4DksjLNr9CzoP2LreiQS6MLtUgbBYPp0HOIMi3SsndmoshOEKnq
tFOcofE1qXN5sweJeoQezyLPsl8njxEyt6MvIzv2zfRWvMCRy46ytKNTA6y08p8h
8UOKMUKt2jrR0W7p3ioP6Cz+oYgNcqbdtmc0a0kFrmPWWZyB0z5UTEsPjnKIbTgG
5lfxm3X3RSl0OfvQv7pA28OW5mjugnjqolBo/K39HrxhIDjyOFeKkKjyOVaiM9lv
MsMOLFjDMXShDbXMFXplWtQmsoHxuaD68y7Kp+XPERG6lU8S2G0WCabteqLSEefZ
58ACQeyX5bB6XCUOdcxClOBEE9wfNqzhwwBcnl9yLKt3DSabCKQ6HevNx11TlRPz
TWE+3QeWGXU+OXXK6xtvpbuixI2qDGymbfiCGHLsOiLcNGZLX8QwXV8pA5O6weuK
YWMocXg0WI0ryASDv30hLbkzla+x1P2GR6c5ccRqyxYpatFDKuuLDSlU8DBbdrJY
jDBp694NJw03t+MyNrC28iTT6WSatRo6wRUtu4lG2esQTDy/KTX9ievklNZKkVDj
5CPq4vJz9W21x7vkXnmLKE8pueiiP7zcp5aKuStpWmcodSQ/ZVNNSx0jYl+Kya4c
KpozPB3WiEUMSN+HdzMzwiaLqyhdUVoo34wnlbNJoP291nsxHiWxVQlg1VJtH8hV
4PLrC6FjvTuMmyzeUJp/YPvPY+qyOzc5vny7H9FoUyA5UMQ46sDTtJrArV6NFxCN
8hk7S+L7jLDR/onxHwDLbMUG4v8jGf1hIwwLRzlLknbO1qm/LWI68dPjklI+98x1
Qxaj5w1lrwP4EbDMtfwltitnZqBpi5RhM+8LX+gzmnHmMeOQ8q3+73WFD5xdbIEe
RKX48SzftPAFcAECBypPm1Acu/iQ6XNLtn5I17K0baeu/m9aTH+/Sl/abYLR/uvc
9m29Ns57p/XKIeirkbNJvc40UmY+6pcdPhm7rxw3rZCDuj+YPmxye8dh2plownRd
RPEFKwErukg0GcsLnhEr6RPRdCQxnOj30YX8kuu90E47HTo3rJ2wOmiYi9bVU3UX
IcFbxQYoP05vWgvR10+IJjpnYKp/X8oDHU9I91HVLjvYLEseCRHOXHh6alHporRI
aLDMas47brfsKWzcP3o2ESdSNzKn7N8SadDsYu1mLopvh12dsbI+DN+ojmj11oJp
r/0Kg5Vd9R/1lp24s8gkuNAkpMz7geX4cgQBaPv7bgDcy2KfAXkm5W6aQTtJbbTX
0z3x8mUEjGBGbAl5xGaBaZjSUvQ72C3OPnkEBKe4ka//cGqGvqrvGLxLBZ64lASa
UHKNgQ6nvOZn5l4c4/lL+35YynSHPqI19w1jy9Q9geZzISLuBjYEfdUwM9sEKShQ
1TduoaxqyVrmxGx2RP6tWjWNbyhJtlMyzRRthDnonU3IdTW6lfWK/7VCvtMdjBre
mSZvhSfZpeaEQoRp+P/dlJDpofgc9vecKC3El3TJIS+dEJzjE/RWm//sCngperIb
eI9C+kXIZtwc/L6Xfy81ArylBvzp28WUVpUozsz+D2zr/kjE5MZm32tfm96jJasx
gIRcFT0yZDYfukPBeY5U/WkvbEZVHsrmztWIgyBIbjxDG8MtQ5T44oNJjhJEbOas
DkwfZdWUBLKKBCzY9KC/47NGEIJ4v1o/GbOStUU73NzQH5WzrXPZakQl7CoNqBlX
F4en8IFfMfdi3LodswjxHstssFk1dePY+oaIwN7AZ6Hd+yRD8FdGp7+JcM3mJfL2
01sCefYsb6Y0m8s6GBgiN5iarrWc3S/z8c0zR6WgVnrWAvmnvsTnKZSJ1VmeBLof
uAIWruIcazpkv3IF753rsyEsT6Y9RE4IJl4eDL8e+IdJrMrUVOlhohD+ROCgwuRC
uwawM8cTHmYXXJ+j3Ytc+U34vL6TzBNP2vlfH3QARtsllQjF5IPEUCt7ml0+yuU1
LZfuFafnOesdnxPayZULbqzlgrTQ+36qX0MmrPvyKiPNmp6Qsd05PprXuC1I7CSi
W5IQcxOKdU6F1rMiE7s1WdN7Gpo4+QQUtvHaOia9qDmj9maudb06ibsnQXvFctSd
734QvjP6cFIDZFqiyMYiEQKNtztaYno8DWglPgJP/Qyf1duL5xreoPZXOH8nnAzU
CxDCmacBfrQQZBq6hO2K7t/U96ePlECwAWA5bwpOHCwHeEGKSvHt/DM1YnArXvey
90tMvCCcXYgR3EgTgJODigWv7vccfuhAV30OiJUTqWdTAAHJR80IKe3KgW0Q6CKn
OWIOSFtTjv3tjYSpFKg8K0LrT8LZ4gotT419pkDka+kiBb9t22GDzqbF8HWxnSTq
vIR6Fyw9gbuQWOOLc4bP6oZhtwyElx2j96Dcbh089DtmRXGDUoqb8CWuTmCWDPYE
fGBEac6Lw4xG1JB1WeoIST9e2hILdVAWDsaM1qJKIHuSMqWXA8T1MGCN8D2rB0Wx
UkE7WOP5Qgi5EM4/cDQWrXSHHjJLiVJEHa+isUmLvDRuYpcld8T438YYwaowBZNR
6Kd1dYcFLnikhxd3u8H30tEIYirJcsr5m+sZy9D3D24OXML4kp9ccDyCCYkzDn6R
8TC+Z+66ALQkvY2D1hm6ueXmoT505i3zp+5MYfAM8FZVaG8LpHzGK+KQdmu/7XoT
Yedlw/kMQCw2GG/0mRhqogvvYruWMZ5oVfmM/8PnSV1rqDIGPjKhkoyaGKPFDgTL
BbanUTuJn7SXNN32oEfbsxr0B0Sz8h60ieP/ablqfcUoQ8WRL5ZFfaZQuCEo7yTN
sECeAhxawHRbsIXI7A5s7SoEl8YSNB959Nj0Zb9sqirygIKgin1fuVUA6FclYia0
96f+laM/9SbgvhNNxH+6Lkv4mrgYZddWFueP/IwogBNGz0+lMb1JShiKvQAHQKkz
zIa5CfW14VSWaWJSN0EAJE4wLKQWZF/a/YE57m9fQ/8c0IdO/lIAksAsyrpK5wad
FLUt0unZkvpik1vbOrfv0QX+7mUbYDIAWr30vG6f2mkZzFbad/74gcdXhYl4gpeW
MuICUaOE8e9OZlZYT3/l5eJ2l5EELnhJBUjlSrfQzQZlVLsXdfA3mdBIjplvNc1r
1+cpBszTKmwjYCCNqHt+N5aRrqVcv9KQMjHT18pvDSJ+cZsEO2YwcbDc0jttyNkG
Oae3+/6+RrpuFQdZIjpG0c9Jo3DHWCHW4h6ReNPd71dbUuUnaNQ8pNfn14A8crly
b3Rhm8VkdjuhYTpuz72pfREoUZciSymLe5yjDnJcgjQ4nHNeoQKLUHLGs1k52NEI
UxD/aD515vFYjHI7rPtrbt8rDlJBWW7MMF7+QFeqPVsZ1Ys0lv53IRoeq94hfzyt
IzaAqgbJTrEm+wNuVTeMYQ68ZdOLlxB43W3plVoHbWoi5QEcoMzHXRRwotdH/GSA
cMnXMK2LXqLyoB7qsPE45sP+by/e0EdWO1v19+nS3Q/DdWDIN7oMUzMoxVfLWDA2
PzHD6ruV2yKQjcMKwlMsWJvgms3lV+0IHJitbj7FsOD/ijCeic1MGLz5wtEYC9Tt
VfkXYvsKbPM8+6dXnr9femRR1iZfpYxBzEKSvVlm1qqpNLHZvPWIpRc8ek4SU7SQ
fwRJ3yLupXWc7Eh9+i9SbT/KtayVI5ERZYjRXbAQNb9G8pOiE70UV6BisWNfkF6s
JPBtnAIN0XQDehVyfHclsVEWi3YEEv55QF2rmXRvxvdL0E/Y8yDDizOZkSgmkh+N
fnm3zJFvTAHGfYevtB8iEZJQaCprfRogJkpRPoUvEfUtXwn/CoeN4We3nNPozvym
Sa90R2M1g0BwQHPFuArJRZKUx/LeN2DRiCt9WhN/mXektj4pB2oCI04m8ubdhvYV
oFpHpVlWDLCJ1VM4WLAXwDxnheetKNUFCnmLooZ3XisaJl0dIXyUL5tRG4tYK4yF
muER/KSFxrpyT9IUoK8PHrSA78OsIjJWJOqbufIlYFhrsNbJLPKHtxK4GHiBYcTB
U8rbWItpWS5/tivVgsBtDG9TfjtP7DSKHoZVrNVgLU5kwfwfYo8Vr0o18qzE+9h5
8IOU+PCAs6Y3G6cV2dpu9YlRBHOclYhpLUZSYz5lktvGtJtkmyDnvrIhpahqaag6
/jNsV6y5ddKNi2R/rd+e2FhZAKUzahLhZkkffyX1/1skg8TfbPXmwKjRTljy7y8N
0zedlzxf3ec6cWBCHhAT1Toohs3ZcWNY45Hn4qo8sTa86YALAe+LXp7t+mCR4FJS
V+5wpX1Oug0Pr+KWi0VSplRBxD5OxDLl8xUP6CeSuSynNvnzRg/AaDTXRWoGWFgh
WRJ+W1OZcW/Eru9FQL3bHKbm+XOQFPT0ODZypxygwLygxRowXyYB7WJYldqVMsQW
kVteOlPT8JyIKfbyLfLnOn3N7pNPFK4/RqiPxyVt1jwougvbdArtbMyt+k/yqNaY
XvhQXjRol8QDJHvGZQIZD3ONXezMsRu5i98QSUvajBtc3G+FXhNvM7aH8DQIJTOH
dXgge79e9QYZ4kaUNA7yYxZnK2Soq7q5jbydnlnJJ46jhKteoZUYuWN1MQhl48D/
hScYMGwg9UXbYmui5DKsJdLUMa07EQkdtK/H0EfYEMfHBajS7gzddp6OOFpYoUCA
3v2Y7KdMGbQOHkUfvrW8R28eCI8pxsWvgmksmO6tgWZOR19gcDIIqGvBFo/z5+04
m+2E2HkGDCuRX0cZeYpQaPBEo7klHf5QIVj+S+3K/BgylV4HAa5z31qP+IAAoUNl
vzWxp81NTmo/eNeZ7fYzbRwbu9utp0+3i9OBVuVj7ambdAeWyoBRuLzgYaGC6jcn
gXSwCTENG/sgtVok+FS2j36D2OVm5IFzBycQlaEcpqF18rBiCHwOGBYJ+QI2awbC
PXDtyldxGgDXHAwM9lCG9tbEJwUjmwBprczJt0qbgapU+4RpoRMz1Va041VetgQG
aXFssQu1o4vXS/dly12+f61iFHxJxQep1/S9a3ONblDBNlVi5x2zIwtZBh9Y6bYC
B59QpZi0XPY8N1gcU+sj3Rbr1bbu0nnWa8c0vPbpTIyPbaD81B5jpS2iNiYmmvHf
Dfbix+p5wBhBa69UXVfCp9xdI3wTYUswh7UjpRPkh+rHde+Fcz/Jg2sV3gaQhLkj
ngSih9b0mWC7JTNATnLNF9rUsG6PcmnssYdkORnWHAJAjgy17mRRmv2WezuTENuL
NGsGKXtbcZts/R1v3GKZ7HQaXo8b36eyohL2ksPcLfK7xgqKb//koORcFcjdoT7x
5s3BEMAFsID4RULlsm7O4R5D7m322RXIC7eCpznqzgT2kQnHIlkM4U0AjYd+sn8S
02e+hyWrKVCQEufdk81mIupKcyMxNe7K8SROdysQbb+f2vPGp9Fkm+69lnXM3etl
Yz371YNqJNc277mWj3Smrh2KMOCSvJMKKazTF5NTV1AOuvw8SVI/MqTiIiYyWRQk
f2mIecOs6HdasVddNVSsIKSMoLo8q1a5tpTTGgvJLWjeUG8AIAAI2csBXyHu5oyg
AW+meGZULl/tL5CFTtopFfFPN7f7LaSTjpvqGXUa5xr8JjWZYTOUewoVaizz1TjY
8PNByQjf9re2BJGORK/6hDPkBhwthuJilYO6OmrA6FB54t2WStkAMaFnVk1MYUn4
JA4Ckm8wyxQT85Oh0bOsYNrrxEpUWX6LchzRl3RvWd8Ibn3kdXoJHz93NJ2eoQ1X
b+oAMCMHHFp2z+EHT7lcEMeIdXJfI3aHLN7mG0irR56djVlqo+OZC+fDCmcvO3AF
kY8carrNjv0b/Oklgcvaupq+eZcxrKhGRILq/ezkdXivK5OaKMxE8qhPu9LPirnV
mQdcrr3YNbg71Q4dHfeXnFo56qRXB+FurYr1k5qeZ3p7i1GqTV1zbVJiQPBL1JCv
XjsYsMrLnwxKrviw/2hWa6QqrxvHvJap9LvGkVDGGM96ATufkhUh42Mej6QkU6hY
c3WzJhrB7IqSAQbC48+UacHjknfJ+Ninb4e4aWr+dZ+u5KcTyx+YXtW3JocwWziQ
L51+FhX4bTxl4nZVJk5A7dfx5Srx9+JhouCMHeGFPL6NUYtL+QlfFxrW0mp19qCX
HYUjE+CGEa/vwMY6YTVxJVWlR6sQvLc4eIhcKvO3M7xfc/bpUNU6b6FRXsR8lDZN
YCh76MmBubKYMFzTiaDjpzlObPkfAmw2D4CCurtF5ERfHVlzH3nGhCHo4FlHZUv6
OwJzM0oz9NMAsHcRBvIG9LtQCW2qlLql6dziODLkQci+Q0ENeAaIeR6WV+SfgG4B
bV1OwOa+QFyTdNc0LUZY29HGp4I19iJtX62++gISbpSZ3KGIlF04Q++V+2DvPkrO
uF+hCqR/LHQfOjo0bnIjMFAo48043yW9v6/FayIk7lYP428iTzcDRWjlLf9MkL/f
S5mXC7XPZYBn9vEZUivC0WjFIwS8fXhyHXfJMdaRQ55TlF8rbJLPEkJd/xCQ/fRS
W9Yd3YNgI1kYn03Wp2MIydTjSSsqX4KFAlG/45mKEFBKT+C+WbgoXGvylNDK5sdx
e3c0XbMcaOInt9z76TgmTTdBPJVH60I7waDckf/l84EgNToqplTRabKVBhrJzJGr
dNXvni6noCzLRjaXl55bfBvrblA9FgOwWOPGVbTNmi3nPLn/mMj4VcE8vqvPWcA/
m5oUbT8TBnoXSXRfP79luzqxF1Xby+Ln07vQrIP4tEUjB5hvzwlwOpzefNii8Tt8
xpQcHTCId6zm/DY0u2WR4c/a6DA/LjgWTPk+5VICyu6X4mGXxnfpTjVzwgj/2Fh0
5i+wprImlomuWg+eEeQGifp/+2xWfNShvSynloUjW5TOpIYBw2jD5Jv62K3M13w+
R3sSgH9dlguzfFzofYxhPrnk5cGlQv9YAUhn7fulJntbcA30GEOyx/+8SiD/0up9
bfrcMrbOvECH6YHH0iWhGCYPjJqAuPFp/1Mi9d8pIxKSN7Ur0nglVtcMG5qyv4Uf
larqCSmdKVzT5LGec9ULmw==
`pragma protect end_protected
