-- wasca.vhd

-- Generated using ACDS version 14.1 186 at 2015.05.28.08:37:08

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity wasca_toplevel is
	port (
		clk_clk                                     : in    std_logic                     := '0';             --                            clk.clk
		external_sdram_controller_wire_addr         : out   std_logic_vector(12 downto 0);                    -- external_sdram_controller_wire.addr
		external_sdram_controller_wire_ba           : out   std_logic_vector(1 downto 0);                                        --                               .ba
		external_sdram_controller_wire_cas_n        : out   std_logic;                                        --                               .cas_n
		external_sdram_controller_wire_cke          : out   std_logic;                                        --                               .cke
		external_sdram_controller_wire_cs_n         : out   std_logic;                                        --                               .cs_n
		external_sdram_controller_wire_dq           : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .dq
		external_sdram_controller_wire_dqm          : out   std_logic_vector(1 downto 0);                     --                               .dqm
		external_sdram_controller_wire_ras_n        : out   std_logic;                                        --                               .ras_n
		external_sdram_controller_wire_we_n         : out   std_logic;                                        --                               .we_n
		pio_0_external_connection_export            : inout std_logic_vector(3 downto 0)  := (others => '0'); --      pio_0_external_connection.export
		reset_reset_n                               : in    std_logic                     := '0';             --                          reset.reset_n
		sd_card_spi_external_MISO                   : in    std_logic                     := '0';             --           sd_card_spi_external.MISO
		sd_card_spi_external_MOSI                   : out   std_logic;                                        --                               .MOSI
		sd_card_spi_external_SCLK                   : out   std_logic;                                        --                               .SCLK
		sd_card_spi_external_SS_n                   : out   std_logic;                                        --                               .SS_n
		sega_saturn_abus_slave_0_abus_address       : in    std_logic_vector(25 downto 16) := (others => '0'); --  sega_saturn_abus_slave_0_abus.address
		sega_saturn_abus_slave_0_abus_mux          : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .data
		sega_saturn_abus_slave_0_abus_chipselect    : in    std_logic_vector(2 downto 0)  := (others => '0'); --                               .chipselect
		sega_saturn_abus_slave_0_abus_read          : in    std_logic                     := '0';             --                               .read
		sega_saturn_abus_slave_0_abus_write         : in    std_logic_vector(1 downto 0)  := (others => '0'); --                               .write
		sega_saturn_abus_slave_0_abus_functioncode  : in    std_logic_vector(1 downto 0)  := (others => '0'); --                               .functioncode
		sega_saturn_abus_slave_0_abus_timing        : in    std_logic_vector(2 downto 0)  := (others => '0'); --                               .timing
		sega_saturn_abus_slave_0_abus_waitrequest   : out   std_logic;                                        --                               .waitrequest
		sega_saturn_abus_slave_0_abus_addressstrobe : in    std_logic                     := '0';             --                               .addressstrobe
		sega_saturn_abus_slave_0_abus_interrupt     : out    std_logic                     := '0';              --                               .interrupt
		sega_saturn_abus_slave_0_abus_muxing	     : out   std_logic_vector(1	 downto 0)  := (others => '0'); --                               .muxing
		sega_saturn_abus_slave_0_abus_direction	  : out   std_logic                     := '0'              --                               .direction
	);
end entity wasca_toplevel;

architecture rtl of wasca_toplevel is


	component wasca is
		port (
			altpll_0_areset_conduit_export              : in    std_logic                     := '0';             --        altpll_0_areset_conduit.export
			altpll_0_locked_conduit_export              : out   std_logic;                                        --        altpll_0_locked_conduit.export
			altpll_0_phasedone_conduit_export           : out   std_logic;                                        --     altpll_0_phasedone_conduit.export
			clk_clk                                     : in    std_logic                     := '0';             --                            clk.clk
			external_sdram_controller_wire_addr         : out   std_logic_vector(12 downto 0);                    -- external_sdram_controller_wire.addr
			external_sdram_controller_wire_ba           : out   std_logic_vector(1 downto 0);                                        --                               .ba
			external_sdram_controller_wire_cas_n        : out   std_logic;                                        --                               .cas_n
			external_sdram_controller_wire_cke          : out   std_logic;                                        --                               .cke
			external_sdram_controller_wire_cs_n         : out   std_logic;                                        --                               .cs_n
			external_sdram_controller_wire_dq           : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .dq
			external_sdram_controller_wire_dqm          : out   std_logic_vector(1 downto 0);                     --                               .dqm
			external_sdram_controller_wire_ras_n        : out   std_logic;                                        --                               .ras_n
			external_sdram_controller_wire_we_n         : out   std_logic;                                        --                               .we_n
			pio_0_external_connection_export            : inout std_logic_vector(3 downto 0)  := (others => '0'); --      pio_0_external_connection.export
			reset_reset_n                               : in    std_logic                     := '0';             --                          reset.reset_n
			sd_card_spi_external_MISO                   : in    std_logic                     := '0';             --           sd_card_spi_external.MISO
			sd_card_spi_external_MOSI                   : out   std_logic;                                        --                               .MOSI
			sd_card_spi_external_SCLK                   : out   std_logic;                                        --                               .SCLK
			sd_card_spi_external_SS_n                   : out   std_logic;                                        --                               .SS_n
			sega_saturn_abus_slave_0_abus_address       : in    std_logic_vector(25 downto 0) := (others => '0'); --  sega_saturn_abus_slave_0_abus.address
			sega_saturn_abus_slave_0_abus_chipselect    : in    std_logic_vector(2 downto 0)  := (others => '0'); --                               .chipselect
			sega_saturn_abus_slave_0_abus_read          : in    std_logic                     := '0';             --                               .read
			sega_saturn_abus_slave_0_abus_write         : in    std_logic_vector(1 downto 0)  := (others => '0'); --                               .write
			sega_saturn_abus_slave_0_abus_functioncode  : in    std_logic_vector(1 downto 0)  := (others => '0'); --                               .functioncode
			sega_saturn_abus_slave_0_abus_timing        : in    std_logic_vector(2 downto 0)  := (others => '0'); --                               .timing
			sega_saturn_abus_slave_0_abus_waitrequest   : out   std_logic;                                        --                               .waitrequest
			sega_saturn_abus_slave_0_abus_addressstrobe : in    std_logic                     := '0';             --                               .addressstrobe
			sega_saturn_abus_slave_0_abus_interrupt     : out    std_logic                     := '0';             --                               .interrupt
			sega_saturn_abus_slave_0_abus_readdata      : out   std_logic_vector(15 downto 0);                    --                               .readdata
			sega_saturn_abus_slave_0_abus_writedata     : in    std_logic_vector(15 downto 0) := (others => '0')  --                               .writedata
		);
	end component;


	--signal altpll_0_areset_conduit_export : std_logic := '0';
	--signal altpll_0_locked_conduit_export : std_logic := '0';
	signal altpll_0_phasedone_conduit_export : std_logic := '0';
	
	signal sega_saturn_abus_slave_0_abus_address_demuxed : std_logic_vector(25 downto 0) := (others => '0');
	signal sega_saturn_abus_slave_0_abus_data_demuxed : std_logic_vector(15 downto 0) := (others => '0');
	
	begin
	
	sega_saturn_abus_slave_0_abus_address_demuxed(25 downto 16) <= sega_saturn_abus_slave_0_abus_address;
	sega_saturn_abus_slave_0_abus_address_demuxed(15 downto 0) <= sega_saturn_abus_slave_0_abus_mux;
	sega_saturn_abus_slave_0_abus_data_demuxed <= sega_saturn_abus_slave_0_abus_mux;
	sega_saturn_abus_slave_0_abus_muxing <= "01";
	sega_saturn_abus_slave_0_abus_direction <= '1';
	
	my_little_wasca : component wasca
		port map (
			altpll_0_areset_conduit_export => open,
			altpll_0_locked_conduit_export => open,
			altpll_0_phasedone_conduit_export => altpll_0_phasedone_conduit_export,
			clk_clk => clk_clk,
			external_sdram_controller_wire_addr => external_sdram_controller_wire_addr,
			external_sdram_controller_wire_ba => external_sdram_controller_wire_ba,
			external_sdram_controller_wire_cas_n => external_sdram_controller_wire_cas_n,
			external_sdram_controller_wire_cke => external_sdram_controller_wire_cke,
			external_sdram_controller_wire_cs_n => external_sdram_controller_wire_cs_n,
			external_sdram_controller_wire_dq => external_sdram_controller_wire_dq,
			external_sdram_controller_wire_dqm => external_sdram_controller_wire_dqm,
			external_sdram_controller_wire_ras_n => external_sdram_controller_wire_ras_n,
			external_sdram_controller_wire_we_n => external_sdram_controller_wire_we_n,
			pio_0_external_connection_export => pio_0_external_connection_export,
			reset_reset_n => '0',
			sd_card_spi_external_MISO => sd_card_spi_external_MISO,
			sd_card_spi_external_MOSI => sd_card_spi_external_MOSI,
			sd_card_spi_external_SCLK => sd_card_spi_external_SCLK,
			sd_card_spi_external_SS_n => sd_card_spi_external_SS_n,
			sega_saturn_abus_slave_0_abus_address => sega_saturn_abus_slave_0_abus_address_demuxed,
			sega_saturn_abus_slave_0_abus_chipselect => sega_saturn_abus_slave_0_abus_chipselect,
			sega_saturn_abus_slave_0_abus_read => sega_saturn_abus_slave_0_abus_read,
			sega_saturn_abus_slave_0_abus_write => sega_saturn_abus_slave_0_abus_write,
			sega_saturn_abus_slave_0_abus_functioncode => sega_saturn_abus_slave_0_abus_functioncode,
			sega_saturn_abus_slave_0_abus_timing => sega_saturn_abus_slave_0_abus_timing,
			sega_saturn_abus_slave_0_abus_waitrequest => sega_saturn_abus_slave_0_abus_waitrequest,
			sega_saturn_abus_slave_0_abus_addressstrobe => sega_saturn_abus_slave_0_abus_addressstrobe,
			sega_saturn_abus_slave_0_abus_interrupt => sega_saturn_abus_slave_0_abus_interrupt,
			sega_saturn_abus_slave_0_abus_writedata => sega_saturn_abus_slave_0_abus_data_demuxed,
			sega_saturn_abus_slave_0_abus_writedata => open
		);

end architecture rtl; -- of wasca_toplevel
