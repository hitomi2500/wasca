// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
snWwHIWXxvh9aBF5zH+khc4GJU4HXmAzQUop/11DmV6LAEC4mD49cmGZJgO1QLNF
a9YoQPMwV1k1g69luo99BxJ4yRBtVkLnwYr/l2kCUYXW+ugwDfVcAvSAJx4FMFZD
UA7GNaO7OwNetjvVSJ2d3yjI7WGfqp8quNMCeDAOxR4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 107728)
Ji27YJQ/jLWxy10cOrTYmnLCqDs0Y25Mh2c0rU3LfOpW8/nlxAXsjQKvdtGVndZT
8BiSQUxXx3HqMtbgr2s20IWAnN3I1ri42xtYc99HwuQvK47FKJwpnrT3I8zmjw3a
rTtWoztRyJ0sK7WkdqDX62x9QmXqaS6xqhCL2fwr917P3zcoDwqD7uj6y0CI4gdp
we1+DCc/QKvbL2WN8Ksn8fxaG4/gleHi+2W+rwCO7DO18MQR8KZk7LWhB1XR3Jax
GI8maAH+oURp2CoZqnKW0QamRD5ZxhFsmcc/NVVVelu1uH1aFFOU5qkyv6cWM//E
w3mrZHhvRHGm+7mA9KIo7V9Hc7B5y2IKeZFJeTEGZtgLU0OpjFKpeWsQlWOUQNhp
peJ1wRITgE2ho3BmHbUcAlFcCsfCLKKqZwZZEf0Nu4y4+ykQGVfBzql/OwY1YFVh
gAITeLccZnFM/KcQ8deFHQ7MqHbcEe54EW7X6gxldszo1Rx7GvgZfdAS36pBw54k
qRulBBVMZ5l+p40dxwKC0kqwAA7+c4/SCOhXnrDZO4gAtbF1tqr1BYbrFj1348zq
oAkwaYCGpdCm3/ya7Hp4Wi+zhw//Zqd8rKCRXeWbIYMkFXD4KWBt5F11Ze65lTqF
GoEB490l09I9fhjFpT40tJPmx0Mm89Z09gsitnRsqSpQfxsLLij+k1bqIPCeQVLE
jamqsOf3EqeAfQyVAwTZv2guk2Zf7G+04hHCKoXyjcBbZyKmgdAuy7UYE0Fpmi4h
KWEj+YBUz2n4dwksDmEWcDY4FoJ8/TlUPjK6gcRwVHtwwIhU31C/sFsxsugvN6TG
jlUfjbaBEAur6z6vjzSi0pUzs4Np/rS8L8Y2eYVcs95Ao4odGRCmMFIyiuPGbixP
Tb506PRCdP3NVQ86ZKmIM6BXKtDfARCWtARgr1yEwaIOqbSIurtXSGmcbGHTi+YX
FEVTV66uOCPhMqfoWGzI8koi9YcbE83T4eaWtDX5Bs0De8MzKnoSv83IG6JmiDIa
Tv8VE4kva0hgTEjEostll8QkJiNTZk6zE80Sga5gSRl6zRwQtyxA/iTOMeo+63Xo
Hj77gpw9RLNmKr+mmB/tk8vAGypitpJ3apvOEUIxDj5R0qhp1ZFBti8XmU0N+y+P
XVeVv8fXTQwSrBWwMJAR8eqcxRhmjQUdq22SPIZAONka6ddcpjyHj/Jf5/kJjorh
TkCogn+e4WZBuQxIFRCcwiTpbj4IMtz3pPYOMCA0O7caT6PIMQzzIfRchUcs4rbJ
UGV6uiR2Mp0k8nWCeUnPRv8FKVDAXhNDOLiYBhpsszvneIQQwwoeDj4l+AA6F3ma
huINdlkgp/Lpiz9zM3Kr090UOl3xKS1ZS3UBLYeoALzdfmMj7n5RA/FboTjkpdHJ
xywtV5KI5XHcQ9gMJRXmxb2F2u2Cqe2HKhakNFw4He/YulWXdFS841clRYgDvGea
4uIJxS9ZTvcW15qrDLimoDQ3H3RhUTNIAyE8ppXlXHUPXA80cy4oUq9HLB9jzOZG
SfGWMyGfpC6ZvxyjAR3OlJV7PpSbAfJEx8Mhlc+ooAkyoBsSDvU+Pdlwb2Klff7c
/pt75yUHGWNoaAqKWP6B3crwo7MD7vElvoT23n9GmHe+K+VTkVgTSLS9n0yntHUl
A9VBOPIIgQv+ZODxEJBeQn6SoE8F2Hn0PskFrE3HKIrIYpEVY1PYEmi2PDwJTQkI
XijxCVhtLcn6xcrftjTAj1SSWI/tb2UpHZu/15nlp+iS38YUl/0nypPMcP5CFpQu
UmAvDIr/YvMlV2224XieTKgZK64UY2biofOOSTUYBLt+lhzL4sOZ46pIpXQMIDeo
EOwyOoetVGuhYxyWZCszoc0WJOXtolFvAWckJXjuViKngfDP++i0pSb4MUhj5iTA
rpPZZ3Hstvra4VdRpzeyB0b4kUUl/K4KZF2wajl2B6+AmFHfDo4VBR6Iz5iZzeYQ
Pb3/03nvyvFWbLqcq1NVCCwUA0To14lZNVpXV1ph52DS3ZRn43ZL+zjgttRALvS4
Ov2eQ1Anelb5UmCMhTpRQTK+pi4sHaITfKf0XOum6T8yO6N6qeeloWVE2v5H7AXv
8wuJ2T5ozXrGo2dYXFMFcdQCzNfYqMhbB2t/6gxVVPm6Bp0z84oqX5GIDgc7L2ua
wVdW1ZkFsAcLmqYjDtigd9GV9j3N0YTwWMfa907Qa8i6CfJhGWAIlsTPW2fcl9tO
zPvNxd8R9Lp69AJS6TAC0atNFT4100BuNWar30X8FlFxFHzF2bjyal/DExMEFOTg
kRZmCZCQm95ZgIyahrq0YG1Ph9px13LUfcmlJHbYtiKb4n4EdPCAQ6bZhKu9mifo
jeRQHHLVkYreX2E+c0EReIn61cgPAUbQDlBRop3SHAcXzFZaCsoZzcgk+pWILVn8
LtBHUUYjDILljVqsizFJJ/BvjaMMzwVGz/ywjhdOlWT194Ot7ypOYjImkgNBNhuf
LxclA5b8id3WDsgvLJkhHu3ydQxhL9psSh46xpL+sCFs3fClI+Q5aBkgxPyk6cug
+OqBJJV6zuZzWrju8fZ3oS+eUl9rBOW0hb93pf+bOG+iFSh+ECyyI9hbx2IHm4Yl
JmNUSWwhzkDzHNlnj1A3i8PVMi8Kl4uAUeXByV+e7JP0850w8C7dOIqxJDKwvQb6
GtscbWx3AO7ap6+a9AdmYFPM4rDbRQX9/jAq1Kjrn8ump0/DeI5TeCKDz10k2pwz
4rl4WAOYufhjzjLqZxogG5flFrIVY/V7ZKHWl1tY5vvHeCKDVJ7YO84InrO2ts5V
q9ngkT9hMlrSdi9qzYOXHahH8h2vBa9OJGox4jt9Hd1Ley00MtaxzqGC8dIatkal
zWHIQU86EyBmXBhDy4gLNn4Se4Omr/TvZcc4qvHEjPDn1rKzi1VMgdFMm/q8N7QJ
KXWgjoKXMWExIb/u45YssOVtfLS4ScPESu8L6Em8sYgpaYNSFKTC6j+lwcRCim4c
NVgTXSiyyIae6ClKsDNzhjloIhbmXvpeDUg0eZk+f1j33jlFaUeY1Ax4XNuNlHI2
LZrWb0zxpp7BBavnwqrz3ghImZq7vEEh8BhKnF5BU7PoLxM3I/ych+PA24gAp6JB
9VoXzTBaAGpNIz7yFAsVkEKVb0WC9zrRmkoRF/kKepSmn0Q2AEtuJ7gJe3f/WjY3
cvQap7Ybjk/ww9hPCyn2HV0TQIBGy1Tz7cmtDZinm0Lipvy+s23dIxb20Jov37Og
Ke4Z81nn7ejyE8KIu76U8RkUrAKWLY9g4ZwVlhOQI5CYxmBRorSS8wdM62D6vuMz
rs/VmFlJJubRGWPbn6n8fcHgeeAu5S6ZHsLCK8o7x0E/x2CJkIQ9Gnf/D2dVwzG1
ks7gx1QsTSppinIlGRU+HJhDmbyz+AV+zUJGIiD7ZbrPQmcOevA06lY1K1SSuXCI
q2sZ4UnLNW8oqLGEmlWAiwqv9V1709gvOsfLo6pSxmKx7bFiDeetlMzPzW9+AhOB
nC7JGUfAXvWp5K5UDCWB1wU8sjeZfhIT/IzlRfD2+Xigy+t/xqkpgg+e/oEK85n2
NH8hDPJhqsKSPyLk+DktckC/N5gjL9/al6DmrbG/13AG0vEA7aIH1EwIVbP0SQ7B
f3urz/MREt0IhFJHoPetrB0h77wGdHNpquUtlARPCzV463zESF02bJ/tX0CQK5P9
l2CIdjzY4jeOt7Hmjx13qykA/uFDztyia3sDLb/p2T9XCC5BXB63Br2qfw27KPT6
5e9u5veItkirbr7mFZvVgggcB70GIkQYx5NLxPI3fFGlKo79ICZXhSq8ZvbNDHQD
SOczQXhDgoWaqgSxNw/FkZL3I3QDx+Um2re4/ig8yTzevgNmbZZdQSjVHzRaDzdr
cg3y5TNomAlnvcZ9wYTLUzgxoMWrPIz+gu5HELV2Z+EerCa7/O+pSYr7K0HC8CKE
W8bzTDrSwDOn67xmaSLQ6NZUuHnXUsv9y76Og1w9yItQ0wr0KP54CqIrsu8X8K9R
XoOBsSGI9btKZpAq901ctqG7XkmcoDxjb2Zzgv0qDWea7clLY6IcNNBlCoVpIjnQ
obtQmeOtyPoHGom1mldqU4y+YPcBD7rDzhVRZJVkGkJSQpthkFKQU24+nHSqokOe
YwllxRWuxbel21/NjpBmzq/jBeX+t5hLrM2bI5UGSgvz758r846McimgJaBy5sN3
a7snJZCtLW7q7heOUa0eOY4ykbnIBfSzIFcCO1II6N95mHx4IwnNnqC4nGeEvu1g
f0qPxBiuq6FVC79470tk+MZtQQ2eglqh5zj/kk/V1mYqED0SguTZwGhZF192wEdP
gUBZ0N7RBBLw3OdgO/GE+6y569Jrq7pUQLOIt3Fm4Lqah4gHHh8cYfAr8/odz2l4
x2B4ER748UNVNZswRfRkOGrMQ8dJgVypLQimO91XAG1/m1wM+gSpb+wJbKq1JFXP
5bbfSmDru12wSdipcwDX0p2wE2kL+Ix/wc6hqgpgPTa16BxP5dvs9qRj4Jf7BqMK
ZiDtHipHBkZxDHlI6/UcTJX9IApnHD59c8ceWTAcii0iGh+mu0iQQC98YIvJykm8
u1hrPSsldVc/g1IwJLyHHKyDPeW0YLqhgEPLKHvxfuamID6vLgeEFX+f4bMJsPSs
C3cwZJxsDRp2MJplMWtW7npKNhxCxzCxfhiWsQPPFlTu6RHoFFApSXkG0vHMIOAe
6fZn49OsByalPzrdNe4/l93UWDNDankRRiYM9cAm5226HRHeRW6ppj7OXf+NWhGn
XAsun0CTAbMrnvaTB8HWT1i3xnEpGR3aP86b0n33rCZGGAtyXi/unqroO2XRc7XD
vVrcEs4T+Qy0O9tN94Eoez/31YL1KzHiQW73VKXIloPUBpJjtZmM+IHcA+7j5smR
NvxnqhDC4Dyrw/wL/DjiT3hcsASfGyg21+eivNFRyZgo6G6SgquEGzcN0fnzq78/
bB0lh2nQ9rwJD1Ewg4gweFVc4ZjQQW3ZzO1BmlPbhQZGNOPuxbNxxbleEsZDi3bf
ELfM4h3nBgV0ZyI55EvBTjDZC4X55Ceh4Jl7PX1MQhgj44AjhPhpollqd1Pgmexb
uHkC4FA0bfRlsh2z6RBHXs1OavfcPe/OLhz01/uH+53rCLbpqctG5Na+3BiXfzxv
YzPkjALBO80KFsf3StRMeEed08w/wrh3UdQwwtnE7cJ94KngeozJNMmoZSxEi0HY
ZrAkHAcQX1WfbpPIUvTuBOPOgg8vBCEvSh1Y+bHniBjPQ5hA/J2PSiZyHIM6Kglk
ViCZFojTF6EKRpzmVOb7SyuotYp3dgcPx5r5SntVEfzUpLhTSrT8qAVN9W81PJIA
2AoT3d96Olqnie/eJWGUmgryU/4AX5g7pYfG+12YPr5DqEss/NncCcbTLrQ9v4ST
ITv+u3i5AUfSqqNQJM1+s9StXA3CrbLksVWsFJ+tTDCxar3SLZhh1ek/ojZmXIG2
lnPRZ7YPqxm6QRZs0mjIxbz2ltgASLLki2raueNZhtx9rdp1nrUm8ywuJQKxWnlO
mxbtFXR55BG3oe2Kgl3FXNt//slMvpRL9I1hxBNkcRd4DBsYWkShrXsGbvMCoEn/
yAncpCb3wNr397r5yLa5uHPDC6LKyZvJiYETW6pgSgdHp6qVkXCbqWkZKGGEacqT
Ik2qkd97Vky/XtwFf+wss4dAQTP98h6nzTJLYUqJ2Ppybc7Pl5UwZ92DweJxUdGN
PggC2Ur04Y3/PO04BIgktEW3llgsXwX2VsqbU/opJZgUsKgxPPGLKAZlM4AFXis+
ekSeA3wRCjbVEZ6m1bEkzVkd/t9bna7z05o/mvR7RUqV4Om0u9OgI7/TgYusFQdE
iAVofTpL/FRTpYq9tAVTZOmv/UACKckuTQ467HRXHnZNHYgRLdeAj0k97sdnMU7f
IlJFbvRdsmNJV9/vWysfJhlIte9T92yn0/u+ijysUjO8GRd1FPIsepATXTLXp5H0
nfxiwYuBRWrWhJGyP6WIu7VjwGGoRrdCbBZuZnUuisLHH+3gu4TZPfRFbuSf8ACp
67NbP2peHfbO0NIL1e3efF6TEC7nCWzPqH+MqI3EFvF149qpI8cbc0PX1/w9Wg8D
IL9nEpUsO+fRb7COoLJKD5Rw/KCUb/98HhMv2+JFvfPBiKdJb96GAuj7k3B4946W
hZ0oSvn+/NgpyGnlYSoMDhZnf7vx3qRTLUkPe7D+4I6NuhsS977LWvUzxJPBhsWp
aJi2lIHsnyl85ZlsPN6Y4lSRwAWidnBOrvR0TrnZIUuiSEbqO+vx9w5zPXJ+kdsT
Z/+jpszGUJLUAntNLsKHT4xDZBkA3KnUVsJ0Pyr8h0okNoIF1IoVmuhz4w8jdC33
cIyxs+MgcVJVBVhWzHjpnR8Uc1cC2pNQiPtlTxULkxGw0+uenQL8rZwN2c7t6HJT
T3AGaX7s9xhA9xKRcne2KhGsS9q5CoVkXnpWUTKSakdTVZvjnYv3u63iRmr/Q9Ia
XNmCRkbpA9GTmS5FlnfNz15QvXA8XPCgd2XsctGLFPt1n5+J2dH5INGYtzwsTCn1
+POwEQVGACLRMYvPQJE6IDmqnQ21GfjREb7sy6z6DTTpvjBn3rUAbgRVH4SEl0sS
Ukqceee3XQJHFAB3m+Th4h+JVbVFeJ0cNSxVQlYyRLE/H08bU408ks+joSWAN6E+
mv4c7yy9KwGL4sb0bcoQEXGiCDSbVKR50CGGYzwL2D1Ajqvbr5h1JhxsAmNGmbG4
0UdLVU43KwyKlGdmDL9pqWo69EP1Hco0WdnR6GYASmWyAjcGmqhEl2gwwPO5d99r
5sQqvjLMhXKnHX04nCVP8IX7DHFgfwnBdOmUOliQU1pgEF6HkC++zVUQJIujkmyZ
6eICWvQ05o/k0XUepDG5Xp/vB+4X2Q7/TynYCLiB/Cm6g0K494RfJXdERt8YAFvZ
zYyZX5Mw9T90NGkrpvCJjrwwa+4g+NNOPZPohhF81xaYsNR9ivFUSdkqbbXO8mPd
+sZqqRM7gZuY2NN9z5630SzVEpQz6Zn6ZGA5CvVnNUnGDMsT3JpqimY5QXexeXld
H62vZxFdIp27Y00q79F0+CtML1FVq+4lqoT21CdMLPJCeE1f16yqwb/F0eFnrH1a
9W1wKIfo50Lg/NtIN2eKR7i6D//stsYBWE27MlTGdT8dN/JfP3qVZ3l0vV2HkJ42
thglsSZXbrkLcW+q8OL7HTiDieAfmJ6RRFIVhkLjU1os5t+i5S6V31XpEvHNxPdk
OdijJDnaAoQg/wS20VbUVKtpZnSFcZ1NxNiy2leCzbXH8K+2fh3xcCyr+1tr4LVU
PKfGCScAed/hiHF/jopQjxv7nskR1Fve+Agycko2H/Yf7nOXtyPFmRpYF+sK6FdE
LhOB2uAuIWkNBxrVlGfHtc3av1ArLZFnk1F1I52NkegDGR3Ccj5l8RXmwoVUTlEO
8z+ig/FPRNyJ7I07Z1EwK9az8DruSoxnsbyH/bffpI30z+8K/jZlhw+MdpjAGxa1
FdmtpBkWtkdg/CTG3CD+s96p+t4Yy5j0ijhnWtBUhRTKPWjTlG19ty0JCMczamS+
Hl5UL40RMX+OzIdnefb8nwRNt7YocbIfyaIrbHWGnXYoZbeLJ/Rzfb3A5otnFpwt
CYUX4z3YhHe5RnvzgFnImX4ewWxa38vbCwTOTDFk3bh0ECZou8+pMMfp+HHrfw0g
hm7JX+sjv6zvj8ojXzyvAbZZDa78gS5NexxARnKjC5Q5TvwQ1IG/G3CMOebkNu02
5FH+ITO33fOWd/nfxzRCYnu/ML+SkHd4iMldJzu8lnMxjGfN4qGECwZYt/GgL6WJ
yQ90zW5M880O3AKVpMGaMs45RhoHKMpmOqQXlmGSO0khnkWP4DNxR7H5JjFdauqu
hkUjI/F5wRZVHRAa+m69YzOIKlWdVLjUFU3GftYDGyX5pPDgcFESrp3BtpfWirsm
F6yKlAvuj5x5BQZx19UAouu3WDXfEMAfWh4MvpygM/+D8oSdZSJvhd5DCyZKu2g1
a6HHHfdE1hziZrQRGdkCkyfLRVCeDoamNbkEYjap9lgz1ki4/L3BgOskKBIpzQEs
M5vr6XBfJpKsYHHAA3eLGCnq0gdFYNG4dbsuy5BkiDme4+152xxmeM718Jqx6jld
yHhezZ/mY+rjBy/1hqNiXLUns3XhbFNU6cQSCYJQdrykC0RPhCgRyUW6HoLZ8dOW
7gVi8o1aaiCOmx16aAUnEaWI1o3tBxl9Xw6Lum7T97XIBAI3SxYw3DJ/ey+Dy/Im
btr8yPZWOCcvkCgumCYcfmTRB8vZ97Eqe1keGf8hH6y7ZOklmT8I06b/exKIgLaR
rgNeXHRCqnx+bmxFDFMow2EiLTzWIxW1nS1AjEabtaP3BaCGW16/UqMhMzcnI1dE
do4bUWnQq3mpo5nUlustfD5wvkbxt1O1BWvvEUqCPKkn8AuTxjB6ZXPrpeVoFLC1
rK7FAT5Ya6OfYhkGsSmyq8aZh1UH7tR/g86roG6pE7gxgqGw9BWFo5eeW8g6aQGw
P05nVpaN++3HhSCwu8j7bRRrujxsHTBGl/OyObakeeQstgxeOJtrsLbPx8vX2qI7
KfL4AYSkqxBXSF29c9O0+husZNgLaox+82OsSKBpDReOeGkOJc/+1kUaYf+EUUbN
QVKqFGDZH2iWzEjxPqmZheGpXy/Y3lRgxvYORq5nunBjcNukKU/+sbswPbCB3RpA
SsA2IGF4LgwRG8p6NS6Ai1f8KDMYS98MoL9kG5iBI55xysxkgnFXUrYj+ZiS60hs
B7MNs9QcUpfdS2geMctTnZdmnWzWE3AWCGX3oo5+KIjbAlelRkUIF7mHDXcs4esZ
X0SuOpS/NjJNdgSgQHnWpSLA9FROUotJVlTiF/ckdTK8WV00Jx+z6atdtTzbCPDl
6NnmN7P1bXPi5xWt1RDX0pbHjx77cchA1lAoH0fA+luwoxyXCN+5BlV2OkNkTCd7
RQukZpoZXfLn1IGI6EMEvtUVN0qb4j2RKK+pfy+3aZqCK5RbbiZMhdLgSHUn1mnU
93VT6ei6ctIQta/df73nTDWuQROMxh0ZrOwt+E5y6EUxHjDGN7XUEVpU+uDZO8dT
n0r1YmwOUQRmeGFf/H0NTQHoEeNK72pkTD0IB1pVvj8nzt96k4l9Dr1xVWM/fDxM
m6IRqUtTbt/U0y4qRvIFP4h5lWiADHiDtDWosK6Iw5dz6pYyFzDE/QS5dTVgATF+
9jG9qBnMB2vVxJ3xIf9NzXic5ZgIjxGiZKCBOeZdXtY5gBSYK9qlv5U8yAaqe81L
+uvRcQaIgKXrggos4SxwCqFLXsHwk3/AGraSblPgR/ttUnYIQZIsFOsXm9SAFHby
swe7GQyPDYoB7bVBewW9mME7yM+Kzd+FlB6okHZAhnv3F6KuYJOzwIJXnGoT0EGX
o/r05v92Z2LFnbiRsDH1ityAnoXbLZikZ5KGIVqTmNi+cLPsBXcRgcqF2ZCRFvBw
4U0RoWPdA2UmAPcTs/OWLsj/109yPPcUQZCKdPGm8KOkrtTCzIKGsP4s9VNktIkP
qKNXEgrzOPBhyWRYG6EDECLgnXuvJOvDD8Oty08tCOK/CnahRdr0j/ou7dzcwB2D
PVSls0mbfGOJ+PYV31QJwwkoCYgvOKK5F813xR6O3oqYRV2avJn/8sc9p6zi7PF5
p1QRujHxwm8c5C5COwybS7l/7ONEMx2r8kYnqANXGF+ePL6U09SuxMsgzuhmXa2e
OgljOoyjvhGRTLNm0tSB1guzxHN2dptzUzdiDC1KbY711vKUClAEssludkiLjhvH
SyuxSttQ8272dzFDKElz8qSvy/qawn6oIWP0nfyspTzGiysLfVVX/i6xgV8e0cR8
wCC+WOsAM05RTRgL5d0J40SaZj838kva4embDSfgWxlqVzFtI/T60UXLG6c7RIie
3OAJg/8FfPLkvyH+iC0SZU6e7RiG6tj73wfS5O6ZxM5yJFl1pC22O+xSYrghK6yF
XEDwGj2uP6MZzhBhiqg4XYO3WIbT3X8I2GAfvdJ0z0wW/xxgnE0zFyTLfMcASesz
wFTQ42AGjYrws6g4qO3EhqABizHqTxmP+EerqF3A+BBCryjeAhuAlRFgIEvCPG+C
r11VZlSKgvtAZEiZYkrhYRroRSyla82LwEVad5cXsYQEgwaiA7+A9dlpvn6YBDrW
k4DZWbmwvgMc8XCIdvvTa8XmmMeyTVM12UPKuL6jSr62l483APcsZEsJ/xZ9Xavq
Ba9AezbjTPPDds74Z5fUNR8oDnZqOw9y3MUCJLZdmZKb3j/5wPYnTqMeNQMx6pCT
3PHUx7Ovq+aE82nek2G4uqg0nOSXXlmolhcl097alH0TRC8hI2f7yz00grNjFPqn
C/wV9fcPkNAWtaiM5ll+GZHyUQXcAQRzjbf5P3uoNNwP3ANE3H1e8QNvtFyzQvXL
eBgF56rY35k85yw1CKksxXkBSQZS+4rhNA+SHYogmHH+JrWgRKQ7QjukNDfd1Vom
0JceHXodSkGUcQ1/kq1avjGKgRBXhk5oX9DspamluMlOF50UKe95Ax9Zeo7frUVu
i60NsQXhKZ4s6VNMsqe6E/KOHhQUtIQ+WfXHZQsH7YEJOMMno3yCbN8MvxZOh3xw
eX08lrX9LlxrBjkuNYoXeEYMkSQvXj69QbzLCjFcpljui98hvoRcO5Uz90A4jAsx
jt2yjb10PAWTHAxD4p/2Qqz7btk33HyndBXEvIogjQTCBwvexPyh8k54p0MhrYBN
0qo6cTzUxGcl677J1CDJ8ll85EbmYuFhKTwzQwLpu9zVNBAQSuZJe2Y2SLGvYsUU
FmrIQhm+HJmmAsiWhuq7foLBvVecigmguP6hlKucLyDkJSQnZCmH0SfzlKz26an6
S8p0XawPW/3m8fgGLbNsHwbWKxaMXOBWUaEx3mXc3l/F9gQxWjJdiN6ZkzxdDM/Z
tlx6Gq5U003dbqW1IRpWWd3gNrs8loa1pruFiFLyM3J6fffTsasp+7fEZUeFlx3+
qbzjQQbARXx9AA6QIrNg8GRsjLnCRS+uuiU0/j9dOVMTRl4cK1qkt4NgRP46iIRs
MeClpWFtB6XrKxYqfg32AyzBYGhSWr+aJ8y04ttQoOT+ejdxJwpRggsj4OOHjOwu
0hmRPDa+8/SkbQ2Tz59AAMMhIyCeF8Xk7Wr1GNo+UhjVNU3bVhUaOVdCKP1sy1zv
2r5IRcUHGixjB3N1JvMt6jO8GB2UDNgdAf6N6YmcSQYvCHjnM6sdLMMpvet4rEEn
W0uJAY5BpZH/nPAmwlBBRCRwqFSvYf5bZdcIqnzCt1Hk+X1dKPVj8/KJVmQmXY9i
rEaPDvwPgr9ZmMKbQibSrbjuPcmvoJOiY29jNqWSdlPNdwOvosjnSiGLUOyowJ0y
/LdXFLV/dHXXXROX+SfqK+BgeOPqMxbwuEXKbIIxa7g82ptIUHTZruflU7VWEs6l
lGePdrqL67KXhao6a6Ur486CjtE+q+N/IbhhwX1cPbtNyHOKBaTwhR2R3AgAqXYQ
hN+EJM1haATABYJOaG55EfT3eQ9vNnAJwuf2BNuLjvak23NUUcv+C8AU8PAUV8qw
vxpfR2CZAMkpqdCF5N8bw38EXtXwHY/dWAm4Xry5NU+xCNMFV7iHQd6OO19Gm9Dx
HsWY06czkYshuJ0EQsABYMmN9H819h9tWnGpqSAGOXTv5hZkWJFY6oe33qvsnrrS
WXHC0Fa6Qn7o5grYNhvjPZ2hVhtVm1FbFrYznAdLT7UKjB52RyZNjPH5dF0JeU4K
1S13fXJ3O1KaGgrNt4IQillsqozndiqSGyFyLyxR4TyJp2lkZfzjL5JKqnz0XPEG
xYw1GVzcNb6R0fU5lcfIRRxf/7oB3tXEIeA0/hzLbVuQSokLdyTcMrSsvnvTtiNE
PRWAJqIB4E3fgOmojDwa6qVRmacWLr2AFNeIYBKgF20snl9gx6ha505opJD03EFe
t4HnxVtbhGmqY0ikM9uFLAsjYLG461VslYHiRNmaAh4J5eX9wfk8cya0Kv+x9kh6
NEpYtxwPiIG9YArLDdV7ZIyPrwkfeP9jxOhOZr2A5/KTgUGjh0ZgQ/YD8WTxDj2P
wfRltUx+Xdwul3S0MdAojATfTdLwTemWre9QUUSWZKj7raEQy8pDCsWo7rMT9tZy
Z8gI2/5M6u/nu55USQMpxkzypZnTDMdq6+0+DJj14DnTwyRir67U36gNUTpoN9DR
HLQvaVLWR1YWIsYAlYgI4k+NNsiuri7NAfJiPDV/LYajx4GOYojIH9w63hS2ieXa
hwSoZ+gOi56hGHhiYgfG27xZiiWlrQSG2plsbR/DJkVfEU6g40O1fLGb3l4oxkkk
9oCEgJIF57I0miwmTx7yhZWPCFOG+L2d9L7FkiVW6VcdP7fIOClFfJ46ot0qucXk
CKwqYU1BpUuwGg8E6Kj9DHwBryTTIjoPbQPXTw7UCgyTExNMx1d+zdbtwUVFK+px
3BbSeqTKGEAztRueKchPG4VFLrAwJTnr7ZteGpSQCx+i8mwDx4iU2XAJXZHCUHsS
j9BRVAT+KkSe6OpfS+WWA58Lf8/jKzTfer3RREK/J0bDOeTH305JWnreKEFlvARI
uJrRpSMLrYpxQnJ9bd4Rl8vGHvlyVH4elCPxReB9rkbKk4lSNVpDx04o7zzKcKh3
PDsaC0WbbQU83GkscAYLH0jYYDPabAVa3UFSfVcOp67NS2KPROtJM5jNwOjZqjYu
ylWY1hZQUfn/HHZiIHb4YQs5oMsDY0QJTTgHEdsGVXkumEQTDtXT2NNfThFVRRMY
9o35oJ6g+3xu6Yew2qkMZin/URRavXW/IQvcvpWGrm3iuQiugHdHbqTuo57c12ZM
5hH20aOYnzBPVQ4XyQGxaXHK4Sn3O8d6r2IOwy25UZTFJSXawgYWFcGD4iAU8Lkq
XhTsGmwPUzQB6c54IQNfniriTlJcLbXSEuUheCK67L/oAX6IM+8fcHb3rvcVqiR4
YrLCKBgRcnRUi5Eq1OyqicRwS8v6SONaLldBlf7rej0YymG18lBqS0N+PvsY5bd4
WHUEDX1YmVE5lx59cgxX16CiHdXZrM79xe8ZfTVaTHzXnaF2AB9mDCTMkWTZSkZi
59d4soYzzaGZtaofiRpK1pKTcEcbMiA1dbvzoy8vndLDz0joWGTCQMnIh8Pm7Nk7
bo3HSlQWcNi1vZnyY4AKNjX50BMqhlvOo2+p+2vB8cyU3rG4hM7Z/951GaFhpr2d
pNhYz1IjwFFVEp0HnrGFI2VHCYIxTDE+iuW6yXZRP16TfT7Jle7aZKaJENXq78gf
TnS98HVBM195scZP3N47HLAN46zcFO5dqOQlDdrQ3RUT71el00pNqQ6vkQGC6jha
ThdZb3eg0KIz5mO6FkJKyeth271sKJofFAvLnUqcHkYoqeRjdNgumiS4AFEJFIJG
fY48WBIxYvd2D7HgUyu6giw42WHpYooYz6Edkf9BxqcVZzFuCyAvi5IKX7xVvRq8
lN2Eyl5WauOkMkRwxa/qLCuGKfFApmfj+3R8m3OjXBsd6cDwkazNATMnurgZQpey
b6Ubs4NFIh1Yqi30U1K3J6SEuhA+xbOYhwJu78HkSF4jsbPfRPVpr42/gZLgRKCT
T9wC85TOSLAdkCAqQsUmWApLmHGVS19qhHbVuPuW8fmyYHcWUngzy+bBcbLppzzD
ZIvQt5YvMDTkbnUHld6vpvomyQpGNpzC/S0B9oTBI3uCjQs2aJrjMkIlgBMeRWuE
/vSP86g/b634FRGgI4Umr7gqoCEPp5+GWgb+OZCqeiu1o4BUyyCVb3GhNmcjWHLh
EYQV1JSqY4YHqXhiP8j5z7V4xqnUj03dEKCvE0dUcy8348KYXDq7kj2CfmFxQ0Vh
DRFuZygCdbpgqvnkljQ1EPhL3RwhW2wxsuL5I2G/m9QnvFKIM/igDuPEJkrDchh9
JOXigmRE6PiC40Wj2cNBrFq01vZElPL0g4CBe4za84W3rIOrDjHSlQg4f05KyLLD
p+JoddZt/gsusPTJrCyljBE4THSRAg0DIjlJzv2r9b2p+SYEDzo7KWeppBVw/k4L
uQ8SXh0LwztPSQTPFvB77k7qLRauRvrJ70hfdJKJZ9kSC9ky6n98VwZLmPyOZI8K
Lx0ukzazP7PMUaeKQm8NGj2WWGfRTgkmTxGmoiUAfNkfhcBz1Hy0/c4Fu4bROYDY
DXGoxq9j88ePDXd86Fi2gqlL6GX6lD6SOyUvqMwJERTZTcOmhTLI4dswcXJvVV5l
j2+aUvLFu0P3BEIaz8sZyB7rE6vH0eE1jBz6Nr8Dpdc0HWCDcV5sQMssi13qV3CU
UQNc5r46qgHKVyjPWLzHNv2BZO6FnVNv6SlHf8OgHPpH1uL3VlPRUkJViK+2xj3g
pM1tA6qwbYiDeGUHHoCKP7qvk04/GlZBzYwbHR2wNw9p6AAqDFF+R04VMvbmdGg5
UQKd96ILGc9RG9e92LDCx6Pq7IvdzL2vguY+4N2RtvGpWWF1mL3HpvREyT96/neO
fHql/Dwg0LdNkOHnkoy6MqwyKVIWIkOe2w5sb8GYkQc7+KYRPM2B1ypYLAUwXD/k
l7l6o0DSV5a5AKUube3JO009H0rmSPOSgbAwujbsIhLIWDQWRzpSQlRvQEWv+O9R
1I8zTB4u3O3WbH2UnArpiKsMHJYrLZL0hedXpTZEJTTkCQSho0BZVtJuWgim9qoq
q6Ol9o/jBOqLX4/+5XMYdkmJR+zKQ6m9+4bXniytnlZ2JYx8jm4HkOR3loDtPiqr
gGVeFV8XkqacGX5ooFt9uVNHqjnofIyggDz+hCi+iXRRTM5kyBTLgRcr7PVPNODf
N+6i7NMmFEgUSmtFUFEn87X7O8tKtYgtD+ky3VUV1TAeTKRKoV6rIEXSsBAPhRwT
qtTA2CBugmkhtAKcZRj8gD7+OxKPvhh+E4nudO2gyvUdwBBZv2duJYxT8Mqgp/4I
Zp/oHNJE+gnkAll4UDIWb9lw7mFGtUHNF0P043+k7wCWyadfRz9GsnGSXPvSis0A
k3cWptvjZJq2DgrSQ4MTixh4xctd1RGq9/+MOKzRiY1n4hcmz+cLa9lqD8cfml6P
xHp4rfiD+02t7FR/Idx9be52+8s3IKrO1zrffB6sZftPADb70or9NyLZ96w7fxr8
qel/v1zfo02lp04tLQN7KS5i6o0XVmxbW6GxV1qF0MmLt88BwxvVk/l8I9Wva1fq
9y4JD/585KrbuNJY+YRcscSaOQS5zJ8/mNzKeVB9zvt34rOsBuqiFu0xzewCB12B
ctUGKP9hv/jF1XHrcu4JYaruEYxJCfCpRwEFhUs0Yh7rMsiu9I160vLHHZWRmtM2
gAs5/foZMu3AE7fgGdFrhc8Ca+gjvBEL8F1/H3uMu6TRbROl0ikKWooG4OJcUlyP
gK73tGN5Ea9S9fhBhm1ZvNYuqnguHuc8gOINehcRBwO+OaerAu9nNw/rdnf3tN0R
sAAl0X1GXIoz18P6RjM5GEuaAQ37/ukrL6bfqaypiqwlJDAYms5Uo2/WE81TPMq8
itTP/K0aNW5RzpHPJKlF/94sUzRCszuRQnlJe96zzFBohSREKutK2K8vtZY8sDab
zOoOLWlo3O1zJxWkmzck0i5Lhe/iIuevzRhLcj0cn8MOQqHpVVtuhgJyASIKwbrD
3xFjFw4tCff1nxFdhKN0qJ//LhyRTSUV/qj3GjzwClHjUoPDagGhBmld3dbctiJ3
+n7bVkjEfXChMit/2xknsEwKmFrYkxMYbTI8QJxrRilbkVP49txHVXrX15n2nwlM
UxQ5CcfayJ0FKIb+Z9oJEgjGVszFz3upKwsL9fC+0TB7kZgM0V3BF5gRWoPAuz05
QG+Y6mbL90PvtrHJQEuvW7BwnyyH8GHz5vKenLS6dGMUo3fohvEYbKiF74FIkt1N
iP5prkZVYM+xyYeURhPOTyrlMS9IlxeuVDSMOcODRvmqX8e/luTNJ05y5Eft3ues
fk3X/e1GJOXDzdo25uKpl9nSqYztqDaO86/LsVRvku1f/Q6MoXqGP3YjIykmUoJg
v8BzQFjFtuOOo7NjUU5kcZ9boNrEh6McY4sfh7rUiHLgSvHulAqZ0nqOYE2KiMkv
d88gdo/38n7lnLiqfEqJe8gDCbtpztDiy32d+AF9fyk3of7KIPXMIfdJZMh5NOU1
iUI+qaCH2btzRYXwjfC4/fVuSNCvIbeDpuZ3A0Qd1SMfc+CBB+Yc4ZiiXn9Iw1G5
sA8YCfU3v0IcIUW1p8kN17moWG6DgVZIpiIdvk5r2c4s07lXxRLw23je4Je5gGN7
tocjQZU7+bm4oNZrda8uiX4Cn5uasL6NQS1oiA5R/08MUkr7c5jvhKrmEu6gJkrD
9C8FS8z/7111m+kHlegH6po4njHKejogmCLPeH+KJnVpsbsP126TcLAXZiI69mzA
gTjT72hxld2B0wpbBq+mdilgx4HOzZsKhLOTsJDKhYTumVjqXF5hA9B/axFfHMMH
zzCmeHQZ2xDLLja5lOSBCBgStOXPJPgyeRH06JN/W2S7/LJISCKu+5UJCzwutMzM
s4KJq1sqHSfvMbtd7GWO6p1heCPjpWppayBO9iYQmM8ubaDrXXHDXCWGlg/iACn2
hhZ9T6moMuExrIbY00kVFQZshOfn0nLTiLPl9VoErfHLK5+HdvmZwtSNb0UaAkAB
MPkgAil0I1toRcAmjxpf6BJmOLfOvVV4jqeYHslILdGJTJaciRNGpxNgu+MlgY4N
/r5v9fwy2IMTRU3Gq1SXTt2IHcT4MemCNkzLcgHlKZ6RmYmBtBWmv2ZgVnmLqzI3
mBWR5sDRWoPyebgO4CEGr/H2yguhmKaOGo+vp+EcJ1S8LaUVNwofhR5bNRlcgDD5
cwynSlur89P0Itozd2vL4KpacSn964OQA5gh/M2/QS5fCh+4WlO0Rn2A42iqn5+3
rV9zp79h5wBX+QTUSbfjAJnhJODdMeZkhMgDM/skhC3Rxc0GSGlxqfJqmMQeTN5A
vVgSZFTa91umOgdjpa0IL/jp2jLYlRgtaxuzzucUchSyq2ClWYmArKubJNJ+rGBZ
BlL6bhRDs4Iswnvwlc7SlQfUV1KMBbtEcKaM42Eb+Kig2a/xJ30k6uaUSbPliREW
AK7SojdficueMRmueNkaPtRr2ZrIJ1f7Tp/U97dohsO6AkP6DPv0pnD9Ne1eVZJn
Z+bLLirkaGtyuMu3mTpFtm86kNFQrCG8rRUIsxF6gDDoN9xLfrVTB3gF3ZlTTYI/
RJ9wkUxFk7kdV0nfMLeicQS465SDCFlihUwp/szKIHdokTucJRACQ34PKOuu38NN
FkGfg6VzRFpTmTffuHrW5KNggJcN7ImYJJYs4f2BK7cI8glGyTMLZwD+x8A58uXp
/SmVopWuD2i6tYXKDeXi3JwuokaBgoSnWRdJDm5J9sgTASIIQn+pS8GpEqrigjma
KHhIlogzxehNk9lpjVD7K22rfJIL4gDZea5m8d1XnKv7UidavH00MiqdhPSN+fkf
inajgqCKhgD6Q2pMReTPYkiWdSw0KlgimQwVJT+jDDGA+G0bw9GVWOO90GeSYkKf
fqjEAcKeRGooPKCx0o/AFKrrjyP2i68tKNekSq4n4bxTPaBxy9yeBhVrD0QCWmjE
/yH7AxkGThrFG74HlNdZmsYkHu/7wHPBOpHW6Lyy3fOx4bDP7OxOLCe997v5SeRz
Gg0bLDKnPwlIGDhkiDs6kgaiiVxRtAOc/xFy90XR4icYO9sNnaZgsaNR/eN/Q74B
j4iyCjfCyYFamOUddsd7SYvDusO5ChIclZweSOPANlPS7+tLc19WmUpr0ij5wHzZ
c7Wr4JDm9Ytww9aaNZLS4WcNJfHYMZi/+9IYMet0JIWxka9Esh9tqzKeGgbX1zg6
Uz7f6JAPpmp5rp8/i04Y/EfB/dqA64WlGFMmGFoAn5TmjO8gCmKBUgz4DQHw+2mc
fRM1ho8GpcS4XIm/SV4iM5moKU7hDkWGDA4y/3HmhwmkgR9ptH+VmhS5LeLKRWvN
+Kci4YzdPfqUjiuH7F1QrioiMeFXUjOP0h3EsJluhf8KDBCxD2reXGWW5xLWlq9K
34ef6VVoKUmAriOERPbRWYKaA+vhAFv7HgwszzIV/uLPPWKmFO4GEy8oGGVzqc7b
7QxMC2fhW9aPUAQc96zeTxgJBTrshqt1JgZhnGD/7g2KnOy1uCRhT+9xx2pR4W43
6P3YNzy0uHl6mQDWgCA661/iJAXgFai64F12tReiZS67W4r0+8COHpSC8EAkvc/Q
0137go5+Wu4L8uCcDHwTtn3UquPYj0g7qQFeYMLqOzfXr1wIkmBk3iWCE4z91XIX
k4RL9G+yovD075w+Jei3ZW2tvnRlqI5JbaKqiSXByAAejsOBbGpDtopRdH41D5sN
vfOC4Yl9hn+3JS7Gdr1FWUzA5JlYCpcaBRXFhdr39mMCV+QgwSmNeLp9XXkYkI88
G5u4SQ3ZpNrFfiIxjzlYTxJfeCfFvgY1U3JQVvnPZDl/NKbiwRHXeqFsPFeml8H/
mgyYvW5Lxk7s2m0Emtkduyk+aBHcGpPuAhYh+t7nbfmOcO83LS/8UM1GC9ZstYoW
n3QURuA1OJVT3K6IsPa+5ycyrA3L6FxyKF3NOsEXviEduCmKeNurCEBZaiOTqPBV
WedSrSDacfvqy9boH9Xpkq50F3KXeT9mhMaTEzVgUfR3x5jWT3N2y+U8FKNMXKKO
tRxC5KPLHNuQ7NPlnf8avOid4c0ctk6PVJtBpmKiaNZ/anLeGP0f3ZSuZGMeunUm
vDSO/wcCFQlGQipcXSFb8biVypLjudb6ZWn8c7ZYnCy7MY8TV9Vn/PikUuzSqzwo
MoW8OoYeG22z2Tgl/VjLbzp2F+u+BmkcnAqMgCf+XW6seBtHaUbiJyUeZDwHki7q
h2oySUs58lrgqZHnTGA/IGd5H8IMR0rsrXkoUtxM75h6mBST3GJfBgRrEEL6hVxl
wTMW/hgPy+IdLjnmum6cq9UV/qb7phS0zTkqwsjNRebdf1tZHYHAwk9zffi7jfrr
+iGeZ5v9FQ9F0hsapbEnU4cct/BIL/J9qUMzZguPEEM3i31fdzf3XeSuEXgFuilh
ZaheTWxlRlQvowEjXZna9T/HDNIwIc0jfAtKf67PtdkLWVN1+4YGOumt+ADo3Nod
M+O0xpebnWAGvANrxNRyWz/txTtmqn+lMbhIbe1IzliIq+0kSFCdygJQNgReN1XM
7Xj9teKdJujT32W6YOxLOhoXV+SRFgzKIPeKOrUbEpv+YbrXqyJoxaVF4G9PVjjD
hN4d6U6RNBwjNxv5WKyonwV/Fzaz3KJNlXnaHd7FEA8HIPYb1q8WOQR8UJHdvZa0
BOrskm+beCircHTDjCCroH8su8gaR3mUQl+sXWEQU0k++B4HhAm2/M3TUXNQk0VN
+ELHalKAEjcI6034UBCnUA1O5t/f3/PiXNMPc8Kix42ODFGmsH+6QYQqq4UMq3cs
a91bR+eK16gMZ+KL/ZK31lcdt5qk5VdkCO3PO1ZPSePcjS7sO8q7IZxibrRCCACN
Z3EIxPFFMDUwYb/99g65cZSYAsYLDQeQxbBMm8awxOLTrR856E0VOwVnH8SoMtIL
mPD/ow7jjUeC71JVYt1P/0nvzdMFHCXbkMUuxFDeVrDqsr7s5gtFZBJpw7rb2ZUJ
dXGL8Ya7AJuh3sVTQst/s7YcOYFSlGf6KztdGQffnTZHiFzrTo4Ru92BW423yg/h
oZ252Ygn3R2JzTVjBkdlfp7DodkdupzyAXoLKWXl+NwSp5CTY1g785X0+aGfrnax
gZCxWi9CE35QluY3sFMMEoVVUbivb7ClMFivbPMT9u/SK3f4bDSMi6yxsF3LC9SZ
ZSctcfMlB/i1xtd/JkqG8cCqORsHkzJx7p1johulyhSJVj1xBha9cfhTdEG3TCoQ
YR9fNaEMifftVfLAkgBie8ZKMivsNWWNqKlOuJGVYzkSjnFrdHuPal5WEQ9gxm8D
1MWtBmB4ECACBGJ6GRf7hS5ACa5E15w+y8w5CkTCOcsj3mVOk3iJw5U0fabgKLzm
kBV9ah5P3EsqdVcimmmrJEW6tcqE7FI1pT1P0AjQbtP1cEIyKN7UV+wTiasju+4K
jnP/dQpQ3xRXowwFwgrgzf+2B7ugkpOv8ilxX8FoOKD+BKSV8OGL/sTgWKBQ96ZH
OCQwu0lXYV00AqMAWIJgv5Tuy03VGLBKzmFQ/b7HM5zqKIaJEbwyN5qWe1tJ9sVt
yzFBqSAO0/XIzPwRHEe1DVlIBJpY7kwL492U6KpeE5EU1BeLZOwwHUZVuo3daViV
TaGYYveekLMo6AD5VKDQTQi9ysSHfAX08qczGlVNWtN0aCqKVqHDGEiS+0E7D+VK
ZqdbAUreVnM1nRA0+4dq+7qrKP/aNg5O1sA+jrgUDKbmKBE1I5XyoURw4eZ+Xgqj
bf4U2W1QsxJ1AQUhNBLCmdlh3Jzai/6Ng371phJYCXyFeHPemVtKKCVeUXxFClL8
czXvASJ15UmbafpC9H7qpqFev1DRdQ/YLpQdbcPb+Rx/6gufQlD7td6HgrESz+CK
DcPa4gih6i7Xtl+QcktN6jMqsRvk4YrX/v6mQMY4kGUtqyk0b8K4qYFz4etSbWOP
IkvK3flJvdgvbdB//T1ZiPnBNX/RY9jGsFcFD1a1vHQGuBWhHV93juAdFf9GaksI
7iucx0uDSGi65c4A3IEBNJyCCwjPtu8dPaufVHuDkGfwTS8tnx7n1R1ybjrqT8vt
OWCqpYrrLsSZMSMX5kQyt3ZA+ZEAPKE+c1/2ysa/G6yJ2ruPcM1W+bZtKSkoXjzp
2PxHTrbqCnI/akfFVNulHmADm8hKEY3mYj7EH7Nv6VTrEz9dLasgJJTlFX4fknik
T3actp7puPKKgusKebPMuUB3/WEn610WrE8zEY0BAzbLQd18im7XpcrKDqgSr2HJ
Ov7EiprzB2KgMUvz31sQ6JeJDpB/Y83vVOyrhOyEx+S2tTSJoZwOXcyorxk1BMth
q3Sd2+1vh7w72dGuM4zoEDtO7Vh1pXB4gp+cEDwsQYkAatf12HrnBPskeqprUiOh
CHwbYpJd/AzGaSl8MN8VYnRv36RuShi90m75UdqiteHY/0vIK4EjbClOrWG5oi2Q
MgdnM8dGY/tWGiERFsozk9SSoKhHQx3LxQOWaoCRspm01LLd5kbjhdMsN3N4G7LE
WtjdrOez3SYkvWN6hn+KlpWbLhuGwJBgkeA+Ewz6S+G40Z+xi6V7Ub79hZi4tO1I
pkMvr3stxjOEndGfnV2+XTvJgJNjjaXTrzmGOgRpETmefx4v1ugM9ZQFfaHEAbfd
5PgbBGZFtNAxZ1PuRXK0WX/KWI+awGIx6yAoNUc4Ur2XIiXYpbLafm9jb39/0EGu
9iTVsp0mNS+U+R9EyhdObt7VpCIjDpgTyVElfzZ9XQ+wVtjgJpaMB/3QfmjssmCB
3L36xynx9qBOyHfU++FjNpEZTSW9kzPVlIQHATCMqjWDyVLhxQ5gA+M/baQuUONz
NCh6SFiqipfbtJSdaG5tIZKaVet60EyIGpzHKSdm1LIRr+9Jw6mnfcvSjkNV0Pnz
3jUGEODPEq4StqrN1FfG2sxxIW65E2fjDhd18Xpv74S0mP+k862n09cMa859/vCr
PZh8Ob7v/A0M5xrRa7FMWojJypTkIV381c/E0xHXyJbZivwp+8avpEskYIk41Zrr
D94pvjnpaXG5Pakkpq5mQE8cPzkckgas9BGm3a5yX0tsJW8XDjIup0UOWtP+B2u5
tjyXsdn17K/XcO+UcNv9ZeeV2cxIVtLDS52hor4UXtsvnnsSXOKDc5RmeaGMicq8
4Oabh1i7hFaGa7Itoe1oqKUxK0foo0GS1hgfWeryeRQftOsuzWpdP4BWS/2YIRcX
E1RqtT45STWAgdeqeJDT9cVGPz+VVv+3LZYeo/fMSIQoiQIZippPj3m7957g7PwC
+KaIfTHDnmOuwHmrewmVZefG4KV6odD2acYXHSb/U43BcfTHkQtUl+ILSi6H5oPw
o/edhPGm57o2Ld+N7pwu3LHjW30hTJr9oftB3V/bc/PkovBt5nJtHTnSyRTgNr6a
DQAbzp4iXy5ePnEUECpxGPz3GQxZxCFU1WVq8/x4q1HohMDIPt4RDvi3BF/XKHss
gqterU9K6u551JFE0Xzfj1qP0/blQi/muTdWASTy5wicTPSE8qpyRk4o9Y3axnAk
0Wdq/9QBiBKOt95V38rpSQIQ/Y4TXowiubVlz8LakQiGNca3LzamNJCP1SBEKaXr
6ciJ8QL4AEO48dUOD0OwOsI2JKoEUu0Ux+Q+pqx2zeGC2JbiR0jrZeGXQsCZ3hHS
rleSBdyYe2Q0sNarLE57qItMBb+cQJfovb6/ptqWmr8rZBOAUUkSWgPtRs13gze2
MotsiSJRcD27VEpPQQYVaCyLQ9ZpuSSiegDgUcSr47aqVilKe+WadUZ8M1jpEsS3
UN5wDgdxWPN12sozOSQX4zSV5YwQ/hixsewbrcE/nay2SLTLgQc2arXd0T0Qs47s
iJmXDFew84AMOdU2MsHchTpz1Qv1jXICP9afO3Da6U+7t2RYlb5QdOqAFH4RHtLt
lTioiPp7Ahmo6NmLEQm/7n35CtMnD6l/86a/AJiK1dsfujXkpiu7igPKbYhW2wQ1
CGzF062u6s35dbhjVjJ+coUwZdet44lmoGdnmkDJXV6WYKYfREt/hADb5QPHW8tK
mEdFRReI8uL5GXWMdNMxFoxP7uC2U7+5WRlr5mXgLllwQb47wXWuJr/0+X/cZ1zj
s/5oE4m1l3uhl0GZ8YlSPwQaIQt1NdEpLXiMoOv+dpJwMimgL7drb3/SEttxfY8w
zV3Gc8MsEJvKlokV5/yujKFMcnSlg9fcZ8xUXBIO1ZiTLNFZma2hahTahrTbWOe+
PkzGy5ApG+soEXYkRS9tNkNEex4B7ZpCVnJPCZ13+OmXpQgEVKGKbVfMCzidxGhA
5DuHatCf/b45iigYmp0/cSjKEFhXlyqs3sNfrxMkb+2rf9nSmKTuthPaWXPqA8sh
4vYa9m1AuSXvp+MncvcYwEjO/wF2Etuh6saDQ2CKNscgY0ltpRXDFTzEUjytIXU3
eOvnJYNPwpGbcY21blvKXp2beIkPlrEXFUgoD73jbmJVq/Yvy21XVF0Ji5J8qIbv
i4tkuyTWqLtZKRojOOdNRyIJwFbByEie+B7/IQOjkLH1E5pd2taAZCNK14kfUf/v
4R35nnARPKyiDEfxpzrMheIe6jatbgGy04GBEbXS6lAlUNXo2Bvhifcx4B1Teurx
djW5zxkYZH7PjrBq8zjHdRF1kr3Yjmn+J48oh/qUOl303K0e8SRMEN6GSmFCLvP6
iV/I39rvtWLWPcupJR/um624wNUZCu28fjYXV/KuDb1FsrIz6yd9pYeERmuWbdCW
Y8MTdPbOPXFyzUgij7+auZK/3dgUawn96dx19KO1S5Wz2ZjE2xhZDZ+CaEbeoCps
c3cFGBehAd5iHtHRR3Q9M0pbc3vocp7OMaXfa8wYuxWgzhjYMcg3oZoxvpbDoEfS
yQXMqI8c4/WMaWy/qVrnxYGI733jIuq4q8ioqobQ1viWAXtjOEDO/c8rHKAwnMib
o1wVSa2vfXFmtHKfb5gww11s8jm7ifP2NPbMJetCYbYoPZFv7+mvycx71NpW7v6C
icVIJJIqkgpg+2qehfBLhkHgA2V0pyuh0LC9VeQf3dYMnNfyD7nMmeUmi8ua7BZj
w4mtOL5tWPApr1Nng+pZ/HRsB77klfuo9+1uu01VIjFzbmCjeq0gsCpPssMXV2sB
A2jHD1Pb9molmN4QaPG7lwlp4ZGSHqY14wP103ZxonLHejW+sM3Er6XmkVDgkPfa
Y3Qnh5pbl9WUJofYWQ/PzA2mF+x5gzP7cKe3FZ4PZRyoKL5FVygccU6unLJZEaKS
yIb/nVYO0uRboTxUS/xp4sdy6kuQD5DoIzDz/QHxia20BOCXVDyXLlPdiMIu08hW
m3FjtNKEUUXD2QL1u6xVDlbiKnqNtXbmINeOFIpVoO2zL3gsrcogWRZbm7GFPTAc
OkvHJRNXwGp0yqJN8A7IwWJG5AqKXHYyWIzd98u2IB32ZJj60dMvpc1jgaTQBRaA
scCjNtaFs30sE69U7XKi19rl5tXAgVkeC7j9KGKR8+Odpkju78ZJ+I7XVdSkTqoO
he/qFRju/7hx1x8v3DvnRBZ+/J9A3s4333YTshA18FOLwyggvj6OdtkMFvNWvOVh
M8qTTdxy3WG7bhLrMlI8XozDCbxT2t20mfA8bT99b4Tz/Alcok/oVdAtyYJ18ZWL
6caUQUvj6aSVQwrVTVOOeNPNrU56+rlfY5rNgOeLOkLnbxMmjDO1o9el1/LVH4E4
AacMfIJdBGuGm1DbdJwVBgRX3NVVakBY9MiOnApcpYf9RAdUUANRZ0ag2Inkin3o
gDDggF5ZYQaCqLbppAggKA8dHi7lVLmOZAUi197M8EKt/s0x3bpdFJb5PHpdxaLe
s6OWopcHoyVLLMbL87HKu94+axNOzrh5xZBzZGMZyEbfeqnZkdCdZ+FyXuIGaC6J
3uVwz6dsUoOBVcfnACTujEeMR5+dLbs7FdZG/7M+q6CoHFzb9jQOPUz03xWu1Pev
NoGvrTD6yGuOKS1XFUk4ldCFvjzjjUEZZxJJV50cOLuT3/XirwVEp2kvfEadmvWp
J+Oxwzcn23s97aSe1/j0UT1kqWAZGhoZLK7+qdUJ/vEmcyn3Jgj1BJrXPMoQqyxY
z8McetNpC6fxW1/0F14NbZr7UPDunps7gVHfZYPOj/Q2zU2ZOPYk1dVFNi52KJ5/
H369hvKIAFBzgiVEKsjokkpjY0kk3s6N7Y9J7QTRDMkwt3vXRlRkUZSuYB1yzPc0
VJkH+b6DJz/pfhTvP+nPEizpNRcvMLT1Wq3AFuE1DDEGZsvRlPuMNp8nmx0XCT8E
H2wHliUtV04R7euvT6VuAJ4tvrxizD/GMG8pKzqCaOuBOjSV6sb2+OA8aLCuLsTt
RCJPZVYeZxdd0UxS7xZ14nlLQ+Ti7RoorzYAS2dscFczTKgCvBNHKOAevCK3O5yd
eNLb40nk/xpFhjgyutQjFewhuyloanTx5u0zHCIF1mzcq6oT9AsgkUN+ednCOtqh
Y/yx+2vl9Q4kcPdYdVhLgzeLTP8mMmQGhEk2Q/JgS3IYD87UKjzNAINkIdr5qwfa
ne8sryRFdDgCh3FDSi0aM1gNn0gKJgUns49/t2UoF2mYXuHjqxquxihxof5xNbDh
2v2/JWzKH2knRPZPMYFxe7vRXjf06Tzo7m1h+dO7l7j5O1pHXftKrAGiibvFCLNB
JIGus0tQSao8opA/pljLuSRMrIxb3oaCl1ROZ8gMnBkad6//jPbZnusRy0fmA0yb
dCMFSoLQFY2TIeF6uflfjQcdu43z6Qj9yW9CpDP0j2flKvPv1HUNYfQhQ3fo2XKr
ymMjNVGB7S8YR2ZKUkTCtNV/jpJ3/KBwNwV4iDBiBizHvFf906phuxQ5KXIJRxgT
biKy4ADKyvr9E9kCVCqLMZ9ZzvqbJUjjdZnCZcEbNqZDOEN+Aqrbdzjp5D74y2NL
OEg5JYGawyWSWcPf19Wv3gy3nuN2M3HtlhaJYBgTwFn8qR8qYwRA/GS8uPHgYfRU
qFBKE6BdwLIcwjjINMYElpCGkzoU/h0WmA51dM31EFqKbS6AT66hcuJFA6dF0PY/
1qAgaBdjSRLKgqelBATBLVxHRy7RFw3mLRuISCcVmYtURSObnnXN28uptXDuywnX
H5TdfK6gbOlV29q2OP20MR/nulHJK/yQb3lUihhhXC/f3p5A7Wx1MWYVdnuRaJsU
6SJOrQLb0+Lu0J6sanDWCrBiBHUc3Zcbq/5SpqsAKmVtc+MECLzS8F+iU63y5058
eCfpOiglkzigBbaAQfbqJPG0WoVbJNKsdsJe0OX9CbhQRiTCQaV2/rgoc3o03uTR
5vtGa8kFWssq5krcCdMoMilrjMelqGCeQ5AwgJOCChCgq3J8+NMpj5s5hJI9nf7B
e4UdPP906xuC8/4ch5L8w+pv0tF7tx43w4mB1INNeZwWyxWtb9aFMQ6/Mmhm9Q68
F+Ll177k2L6vmst+NHlItd935dbaF5XX42bsdHP8vGmqgIqLhYb0DrpjdatEzpwo
2s5NPYFpCwGpqwsbA7gDZ75S/gnadHcdR28q/0VP4rX4ErC41It4QVNinefRhIdk
UpK1xPssHjzH5wPzDaPU9y1msCeGHgzdmMgf6AlGcsj9Es/UyLX0/Fd52imMUCf5
DneBFvIyM7RD22eDMd/7nHraMSMA63QySiMIpIns8+pKCDVHmv77SeabcH26pN3y
PPSyGvEdkmj1EoDUKhsK3fGDUZXj8vtZypdReCBvoUyf1qM6jsw/+v8GgTRTP9TF
CoNEN5w3dMpCMCZf+6Ql/SGX/JjIYP/R5DVTC7ePsST9StqJTzpN7oqaKf19U93L
I2knA9KQuEQFOzrxAe7tfq84mcDzFmj1/+AtdRPwg2FF1ODczp7owO8I4MX3hE2w
DprR2jBT4qfzpZVCzzr/U51zPUuCX3cnlDIQFLsNqf+BZuOJlBIMAf2bwDtJ2Us5
EhsJHYLzfWr6e1D3lDUjAhdx+fBOA1AnXNPt/RGUSnhhwpOAjZhC+cONPNBdDMrY
Cj6Mt1f1PpxgQQQFJU5jD1G7IhG+v5QdBMIDVQmIRJcWxmP9sYZI6zjJ5eH5B1JF
UM7wVoOINq6nqYLE0Cj/dLsscIP1z/Vxd0QUMD3BaRlQhNEfuBV0VkNgfbV53+4B
Qbo4clZwpn0m8E1f2exdVGzWABPyT8K4yXiAEZ3k1asgjfzh/Zwf5XtdWbGYcvv9
aMBdXY/Fg29z3pH9tv7LEBnqHROmiPMCnYj+mtBZfWtICsjdOmjwaai14vQGYfjh
ACl+A+lOoHR4KAK6wpmHHuIceUh1OpXPSaodh/tk9Uy1isXTC9DHql/I7w76IjGy
0T/6c3k3J9zUTKLCfRRyrXfcQ2MvM3fF8cwTJN4RrnhKWkV09PnO2e7PIkzyB0td
FLMc3Nesop0rPOC5GZ1HafT5Q00Vdl1DZ08KNw4p66xD/Pt3aq/quXvglJYbftbw
roiP93W2CSdaT7F3snrUvTlgN8W7ssl2jtk0Vj/DiZe+tACikvqs3hE2grxlxxax
HgPuWaA8QL9xFYi+s1+B8vdtir2RKX/yYsQ/YWRqcnMgtFsTo61LRgsmcIEDuHed
XuGvRlj/SMSKX2TX8NBAQ+UTPjLSsIEX8ZXV6EwlUG0TWqez5CkJ51xzFDwyI4O7
NkAxJmeeEoQLNDUX5DSorDT2T3gZAK8WTBl9Lk4rndVhcRnFSFK2YajWNx+h/UOx
1NzNTHE+iw6gza1RWTYyMORvh651op2x3aR/+cfENfv+9x6136+CAasH9XSFvBr7
ss6lL8k8ij5aZkwv2i/1nt0bCylng2XufiT/seco85TapkYCTh6Ja/GpokNOEqaO
L/O0FgpwImQb+y9tvB1yiIEJb95fvZE52AzRyI7NGVab2ZqWxKNRBAACZVyPCFu3
yYtd9yDttjMDJA27JVdMl80L9mNUuBOjiVrB3lx5j+365SG3R9eZMEQz2aTzCus/
AsT568ohc5t7fWR6iofYBxAmG0SVbiTmaxOwyW2sM/p7WdVs75GCqpRhXpqje8Nf
iqf/iiIyM9z1ZN9vtv1p/8X7aS9e73fABPXWQdBHlL1eNZmPFCVl7vQGOj+56eRW
3cPdgzlCHTByWPyyq5qEvJ0zJMnDEoermsJ+Fflu+sFltxCMo4W8lj+z9aA+8bNF
18QCQqS/4km6WXoBX4b3Ei+DTfUtIMtoc4jrXvClIkBkTb381SWWuKCyut51H6Vq
ccNcB/+5HGyzlfvQoXYHVrn7ofsMCkE/ynuOtfFOurrooEQ58PFucEYC0+rjbn1G
Ol8Sjvz6xixxgBtdQpPaf9gWkdzDB61kiJ+e7c6CH3BVDvxl2/fPLPYaqm2hUhQx
W2WKvjzMHnyu6oNMKQMMUMqirk5oNQ2MvO/8SrlR/3c2dD4tlmtOsSU81Syrte+q
eSE/6vmsUDWYP8S7oahgHer30B9NuTQ5gJNyFNf+J/ez+nTTvIQ3tmgPYi9AuM3c
4KAa1Pzh/7lDLD1t4hCl66vD+sg5FOZTGTGEUHorLF8u+zDnjMQAPl/xgpD58WYa
8J6pERneQaN2TTITjhDq5gQzrm0etULtkktQJfUFUaKn1OIrL+MRN7xrHyMeTejn
m9ipEjQFEJk4AUSZ2vBFAynxAihgDCm/9Yje0MpVQSnczM/+V/SoFymjpbJKcCe9
URR6FZfo4hUkEln9tXua+gA+051pZE0VWIkCSAsD3dBwv9RMdQCaCvJutf7u4A8K
+oIvNCR6srsX58rLbq5M99chpznTlns3857aw1AnQ/glOGpYRBYFJDQqQ+VZKitj
Pf36N1Dc5PW68IU6domGdB0oI43x+NiWDQqkXh2ecC4J1roecGo0tW9CEyPSRAqw
VUQ9/BOO6ZUP79tm00oh74mYBCxciC1Y1EghfYdhRBEwPvYq8JALratYJaOZOsXG
WCJ3WZyj7EdqWy6/nnATsft+lcJ7JBqbw2927YC4nwTTUpijsxVbTI7AnSLOi8ri
1YCgho+glahUGwIOEUFhcDc6OyAM54cR6HV3mne6vYqyETkfIN8IiVhhv0zZ7lx+
tb5wvbi6T2w6FYLsHmM6xfVbvoO45m87AYV9M60Gvp9mNroScmXYVqxRH5AXbnTc
VDrHx7+LNAPNNyUco9Zp8W6Gn6VYzX4G4nX7imJ5mpEcIWrrQ0beX/kvto3FwhsO
mKYWUWjXG9hC7NB5V8FA6IUvSqVO/GSZ2nE9gI9/Ljq2M3vj3EU5+uDV5YfLJptC
XiaUsWd93fjpLhSmH6a5GDqtkPTJKjNiGwD3MotxiwEu+270WvOiLoaHj/Zdul5Y
eB1qyb2I5lwIbY4GcOjD3/r3NiTzFle/WKzwaRwromlzuSzrowZNhGXxZ9pYO+EH
5QD7yIgOHHTFLIhnAeXPXixiZ8hP8YUBa1/hsSBBHLcZ7cHMqbGzm2vrOWoGA+a/
6NzD8NKhXB/453FObUTruETa6dHqEoMFwCD4sJ7QNLB0ngbdwOXva+0UESNNg0pq
GLzHS8NvZ1dpzaHVsb0FlmGbX5iB5tnCxhM4D1yoWKOo+GB25GwP7kG/Hfj7G9Yv
8PysQuyz5MJmvAQh4IuziMDKV4NzQA1vZkA9ur29MSX49IKJ3VLSD2pA0saKja7a
1jQ68uZ+pUPsf8imufa/gO/+rVdWP6Aqrsn/TXSsTChjGwt/+RhbpQSFlmaoazDT
PARHF0OQOJLEIlYcbS6Yc+qU82Kxp2eRjQSHMJyDLhiKlz9dD4cN0SpX5vMZIIMq
EECAV8GtrzvBT7QjGKaVeW0OVH++zfnQyKp43S2F9fNSu4XAV1DejI+2gjOIqUhp
wo4RHERRV3/F79f59JrND7UVpjD4rKF4NmYsukLO7oOJnhAXa4/3JEuGBn/bPxHQ
/X1qu87SUG1bp/ePa4vw9TG/c3/dQPueQIs8vTPDGNYjlfSraLVtva1TXbW0gC5N
JgXjr2uUfh4lfbjFDlZEEp71+n+491ybCpBfBjrrXmiSwlNor/2IQgoDTrXF46nt
EnWy0P6tZqFQlEtSQrVWUx0+Gb3owCKa2nqEfSd83wdHpk4/RF9Zfm+y48GTmLhq
Q4ClQ7b0DN77IgiN7+DNq/XRntvSWVddqm9ihxe/a2dOCqIXfTCxnHnDWOqv5Ai+
35A2WAwC0IzUGZTbEWzjir8U/XdNIE4mwYT61k6DK+9yCEw+PKxY7dt5hw9NKZtl
xKJEz1jF9Pcp7yNz8ZULl7lWWlEkbcu/xCKrWw+QhNFBg2oHjYpY3gutioOQODRH
yW/JFh4GW4vQCPscuHGeWyAxSLhJq/UJhbcg05W7aLly6WJHhElNQrkK9yvdaLcH
Qg1v1ixpTkb6ucQBLKdlCPi19rtxQPndomKrX56wRIVWhx7Oguz+lrMxRooF6LRi
qQitN3ENUZCTWwaylEaYro/AFVBFaOw6+n9yaCYpVQKgfyTdFtSCBcXVO+t69vQy
HxuqflldPmFjbfdJuT66/4KQQguMoYOi/UO37gmCu5sBbECx/EfmJA3BAg4+pTfC
29HcXaMbNlo2JlRBkJasCPo2L18JZsRhjOr+KmZdqZsmI9f+eceCwXtrwLZKitWq
RRMYq3pkliWZVndwkGzGNmdeE3LrA09qRUilpeTm5iOrYw5Mk5n+Z+yqnWdtqkNv
GniZbjcpImwcQLeDR2tepgAEjOZ/6k3TZuomVNw1Rz+OzkXbEspbODki96306nb7
U5FEnckwYVPg0XeoaF1YnzkA2Uy4gViIOHUGtJLhHcqBH7N//tixmiL9Ey5xwVnN
u1iwUiCQB4m08JLBbOunjvYM7hkQxD9cGkrT1ns2DyxatpUscyA8zIWoJZTC3Fpq
simqFNPthq6O11B4yeU/bJH1M4oy5+zacvrG7/gGhoBYq+JCimh9elactqe9HcJO
oLDcGOLuA0r9VnaX7uQJ8csmgTqBjYdr8zZMyB4Nc40CxJnP4QZ/VRQJGZIEXjgR
TdfyYcIH3YtcFisq3Dhs8dzI+yWI/GnGxSCCxWOAwbl31OMDxcbi8EVhmm5fVs7K
gJBy8GQ+sbGqiSz1n71MeI8gIVvhAm4ARdWIcCbPUt9jvxMN/gk6WWn2Vybqc0Dz
G5jFD/CVTL5C/SRmmu+DGwkSjeEE2xSUxGdfMwCUXkEcOutfAhlAlcJ4koEPQ9Mt
aZ4EJtAUMm/K26Jr2F7uNVATu3P/AibEFHEznrE+Pz5hkhiB7Wnyp8M+i80KP5HS
WSr8Hr6Gh6MVP3FRzYbDjWkL+R9z5Ph00wAIhir8/gBdyDDGa+hC1qyDyTl0u3DR
tYrKPxRdxSY2azHmxbxS5835KKjiIZ8xQYg80/XvxkH3qvsRhgwrUffDMQAFJyUi
4uEZ2s1RJl591yKNRShJw3pnmd4Bt7nKqy0QNGt8LAdacH46t6a7a0HsX3OiOCT8
pKazr6YPJvlt8wWzf409E80r87CmWQKqglV/jhQ7zlyzLfBYlMO6jgzDpqc6rM1B
YEcQNO656wr1OCJSKBKeEM6K+QZ7fywtWuHbev3Adea7OcP7dsVecZfgBARnNEIZ
LTWguopfoRDcRrSsDCsarcvHPjZ69quBtMzCFK6Sbi6nB7uCa6CKnRyCvfzdhdcZ
VW98uUyTOEn6KenbUIA+OBUHgFPxZMK1npaRCyhi4IAHLsrVAzcDNZsSjy+0Hx+M
+dD0jgpBWQcvJ8Z83JYmr7+SADQN5MEcSkO8CEz4DGjUYEIp5LlK8HzniG0mgSrh
7vKmaHnPlGi7Qb9eqjcQZihgBqM7TrkbsG6L7Xa/vAiUk07rjwkbo+CCVolA1IsI
GyhDdn5wafrkRCLJo2wVhhyWcsVWSEcZ7FxMv25bPbhSig8UHiv2lmNNufzJIC6/
J7dZ3OsBtZkyKtWf7Eo7JeHtUrKXYftk2cDQclt8Ag/3CzcclVbVNU4D0uBwYfJl
i/955huDQBpkXdNma6KLNQShoSV+ouu1YKV9GyNhmVFewk+bi3+uMYnhnIojrIMi
0eJZ0XiSKMJ2I/WfwMtx9V7m/tsJJ/7TfLd+mwzfK+xSe3RHp85YKNKbKCGbuACO
AjMmRDh/bjhKRjC6wPpThk4S9IWt+J7Mvzboj86rm4w7dXmddFGVHCA6a50Q7jN3
MrAYzOtESA32NiWbjJgrgR/c6IU3MBK8IbKdGI52oV+EVIggdvnIkv685xM5PX8p
CHfvcU8AS97+SL5OL0eZch/7+FKwXc9CpIIAO/9RH8A1eQCpfm+WafhN6eToVk4I
DIQERgrFezfwy5qLDD/9Ewi3BLdUcZMKqAcE9UrJvk2qkU06kOo4ZX8qeKqgNWS0
fkxE8dMZjjgelU4EFmsKux4vybPCNH+YvShxbaZpTHwEr5BtMn9spwOL2rIUjSsa
dyGEoKcPGihZ6OX04Hjiwpr0mWTqzEMrrWV22zPZ5atbRy34YstqIVXpIkm358EX
41Exkz/hH1wcCm37pH2ktqVgz0sBUNX8R4HZOEfqJM7PCTvR13OzoZzfkm7Zm/KD
pv38m1lFqXXOVEgte0V2le2dbpwpB7WH6zp1bSFDUU96pZqPGJW3cBzQWA+Iv+4P
3G8nF4hywYAft4TQU+01hjMqq0LCaI1vp6W6RzXsul8tmvIOpXJgpzpfYkYy+4oz
xxdoX75Qcrofig001rRaPDjoZiyoUrOqCzLORwHPn7z0VTKQUkSzxhqVShZB8BJT
RSpNh5FFwnDlohMRSWteAapirA9PhgCpcQ4qZWeFfl7QjVN7Yr9KpA6Az45EU83Z
hKCGFGM7kHMJ9y1Fm/tJ4VJxm1j0rvN6/d6Gd5+7mfW5cS5U9e1A4FBUyraizh+T
AN4vJUY4HQlGcnrpr8Ay+lYSGmmjJtIm9ckCmtE0t7u0LPmo3uxErVj/zHl63rs6
28mR1Ql5H8ALUFxX860YUY2ys1AGYc0fXiIIGNpP+H40iTdIjvPLJheJNdj2B0dE
Mae4kdtXIQFNHeWbUfl+5H9u0+aJYX4ZJPr7H8M7+r+polw24vH7u8OJtD9dhDRS
d7DBVulq+GTf83lVwmfQPhdw/u2ll6gVN0wYWFOOUklit+6ODsAYrQObdA+8ex7W
rUhoieGB3zll+Z02O7SccYtTWnmsdk7IyV65p4uNZv4L44zvOxXCnh45O3vDPdmU
ecsH012DPLe0KE+va4hg1Fm7U2nczVQF5wxeskQGEY2yJs8iJKsDOn9T/X31fvCb
fUxXtjsiIVZx3vNrzDgJBCJIMlvVtnkYZNJj9cUeNLsJq0o8HAfP8cekYVePvbhT
A/4pXcFCIFEHa9+KNgUHYE7/JzprnMAhsdduuDfwAvnhSInPZ2G15sbH3qJ7m7QV
pRyavLKXKBIDkFGd7rmSoAfxLjGlay0fPYr7vtdcjVKKpzNFs4NteZUTeV1SQ635
DxxwtJ4GW/g3DKnVa7v9pl+I+r5Zquyu8gcnEgoDwrQG7xKDLQ1CbmGKfwYPRtgz
3l1Xfu7iAZKyl0W0gQt7XdM0DR1qHrahHVHvLZA6Mh1faI5PICObUmp02xiKWZ97
6meP/epwM4mMb5rYUMaspkrMkJaQZliEx39d331WYpP9Pq7PoBDLzoGneL8tiYxL
rMDHah81kT1Tw0nUZU+pB7nuhORE6S5/leAwGlYSOrtYNc8iklS+Ilfo/XXMuofN
RLlgJKgAV458gTEw607mP7UucENk8TxzJHohgy0kKN9jWP0DZ6X8kbX1JlhReYiP
rPwfbBWLmODXZSK+TkliEjEu/0s+ZR0EQ/cFF0z+7XgNDjBgQYOMd3KfBxu5kvBH
XhBpt7WY3nVKGA6PF8e6cB23k4d/YvyPNHd542vsv7vSvQ2qYN6U4oLE4Dtyg3m9
E0zys9m0MhpaIUoBchjUCAdb1Wix76/EzgNJn+MO9dGOQ3g564wPihYdfT/sVPHP
9eu4vcR1TtgK0jo2LOXJsFe0bkXhuU3CC3yWDdCi0xiOxR5Jp/NEbYvPouseB5Bt
FyM6Cvz/k2AwCzOXMbskAGViRgCa052JIIKSQllUaW5M82LCTWiX19aeeY9rGKbv
7QabrpP/Xq9dLnnMcuIVhoLhYHKppOFtg+bCXT2Qd48C/njUNsA1VqukoWLwa7CU
oClLnDYfmGDRErrpfs+fCEaPtTrD1DdS/PM1JGbB+hG1B0izN2NJZZ6jrJxptXqO
wV2esFFNWOncYzuToksrkmerf20aCJGeH41zQsuvGz74f+p2i9oMdmqOBFbmECwj
wElh+QCdQftojY7Ki/1/lJSSgmI2sn+/NckFMg7YCWCciEK/nH/gf7PSsV+2aMKf
wzAk83ErrYKKgdw4XE04m6RTAjNEcMRKeaE2MqUvLkjBaIZsuVsTmf6wtH3s7a+J
YtxO/V0g0Qxm1tzLfyy0VWhTxVOJTZozrdpVecbscfqaBLzxU//qn7by8HiAV7FI
aqdE3StzpISRq7zCJRKxUiB6JJbnHN3bRJPG1QdKp698c/mAvsatiP90WvlF5t5z
S2K5S0gmf0AAaTbAZM4DyK5z84zcwwUR6OPnop0NGHE4vS3zfwQV4sR2bZAOSJLY
LVhBqcACBFshZm9O7QkbpeDu7CigC7LQl7in43h8x5yxr6avC3srGRR2QxZmWxYe
Ns6sqBswGx0fNNfb3bDROOjSWZLnPRuVzYuDHvpP0Q9UHMtFPRaR/qzZBph0lqUD
3yTER5jAzsLZpMXa0rH47PrcTYaZA1kOUUziiCx1gHxX3JE248uDx15DUDkP2A7+
qfQxkxF0AFleLe4gYykgUPv9P1rqyHjlhMO865+N+CQkY56llVXlmCxL6NseHrHA
R9Y5Hxh/pfxRW+K/Tws0z1n66K/Bvv8Ts1Rq0Rgkos2Kta7Akh6p23rrESQmvnjO
3WobKHIz6NGjTE0M6wrFjap2mCDn7O2zYY0/h3O7OJzmzuw40NIuHwpHO9P9YHm8
lzI1gcxhxSx7mW7wlox22r1nDFq1DpQ6eRfvCJ6BS9f5fpYDxhzsuBDeA8OYasnh
K7ipOUHkgrNCB3MJHDXkLYIPpkE+WFVVObJla0fUOZJeq75qLq7dwTl/+UT3b0WG
kHPnh0uIB3ZZDDJxNEbWLm1KPbhOCd4EHzj3tVy+2wftwEPpik8EWTQUnjRdN3z2
2Jkdk1eRrf1x5wVrcKN8NpK7uBTpghxEpflEP0DTz2mKM8vg2IjAmPvb1hwH++q5
INHEmiT2IMS8U4WZDqo5yHrn76PLMwgJnABq/I7MXcovHhRrpfl1EOWgiX33MHvz
1jKzYRRWlquwS4coxNmcBzmGaW6/QkU/MWcsmO50idKMIFFwsK1EIiG3oq1CdbAS
tRDDnZh9WlDwgMdeuHpxrOU1bw8TrNGh44X40GJZH9JuKw5GOgDtLY4ObqiDkZtN
6vAx94nUzasNPyppR3pAKblzBhGfFD6jjae9TjsYAqr/y8O2jNItuvniDPHUY5cD
RrJL+LKcXHu87cnDFHZJaRiftMhzcP7QR6zN3mGTyjQaLWfg3Ykudm2GXVep1kbS
KPSxwjJ8/d2RagK4YLxquyqXbphr9KmNqB42BSfKC80Z3UJECakXQ+4d4TvXa/da
YO+Z0SXTs5eMAvrkuzz4p4EpK+wKn2+fITD8MyUTcrtjnzkYERmbcBkO9dy9M3Qb
Ovmm8QFzdBbj+SEZaTDsD7AUL99edIXHVFj4myKAOQ0LoI8I7y9ES0M9UakqYspS
3aBvMs+dE4ITdCk3rpNwxS5zUPnAn+0xTOAZMwgAg0m++55ndu7nGFO3S/IQMdvQ
PKIhLxQBvokNwBaNvzhH20ED01mgDMW452pztE/YuVnD0WeAhpCV4Xmzy3KEYZr7
FT7Sz+zyPP/5Uhd3aiUZnYbYpaDgVnyFavtFi/reVDQn7kruuQfENPXIL3pDDRt/
0Ekp8ELrGUEAC7N6LWTQO7b0dRx7tdQGkMngVGjPsWIkJ4ZnabQ67tafy5/JLqpP
1pbObuKTHFYEB9HRY8zUujAhkD/RhiMVMDL+EIEsMjOFNOh0u7s8NAdE5eGO6wyx
Jj7l7h+TreSxlVxae+tR/IlPm6K1Nate8lkVvJTxXwgSHeSc+876sgca0ANF6d+8
lbqB8FLzhITx1EOs1do/CE9kw1UC88+tCC1nvaDihKUd3eiT1eDJlDnrVuDhGrxm
PrBaAT4EMLTozMQMzMtz382tBT6T4filhio/8LzWPRCP5I0REUepElKaoVlzXf64
7jOJHmkyB7v1RgtZC44dKPe56bkQyqWuMDJtz70ewwnVziVfsZ5QGOKaphrhIrYn
NEHOnnO4Favqv8dPetWIU2Fuf7r5KU7gdF/AmmGZyPGApY9qIxUNySM8avqVHmaf
6+TjloUZNxOaSN3SQSEfz82S4KIhXR4GrmUI99JtM07/nTCEcb96jS4rw0X5/ZJh
T646QhUzaOnpwwr+6sw/lx2WMKQBl+tvJICGpo0WnlrRF//Unodpe5KgBLbnZDbM
Tsf+ZRQE8Fb8y+2qukb/2WHIgjmYk5jGizCiCcaJmWvcQsZiCB2IfWjiYGqj/rHx
hvNdHqmsaP0kyNqjcjmU9NK3W2pkb8RlK5BK8paqMa+CtTxJbU2fO+GjopcNU2s2
19SOWLlQo4DSkExRtX8q+cxA3LzwaML4R++jh06mRF03CX9K4rF/63013LjltMUE
fHr+76717syQ2BLzYO2M4mFgB9mXyCwEI8Yno0tXqmXIvyDnbLINdpnzr0ryVdC7
8U9UisjCqX1XgdsEi2/KoLXekOpWFqDmcvdIsd0Oe2P3JbXFwY17K4kKsHb9R8D8
Ra2Z7orfGAtbGolH/UxCvD0dRoKxkWQyN8iec9vY6tDZhqXTdpm8nPKwxi0PKeeA
LZsULiLZZtfh9J0AxQ1Q6q5jqjkBvc4qwGp+KfbfzolW/9aKgUhn8+TkhpClSPTn
5NS43u6aDx/bBHAOm/SwCVLo9X1mOIukyCp55sFc1uufcGeVg7TlGF3L+NAsNrSv
j6kY5jeFSdKMfSbD4vkZD2GZ8bhvGQOkZWrWUI4IRPI9Bq0DyN60lM7h1hIc3WP/
SGSIS69kNi2F/paZFpMV5s3iQ3hpS3X9ea5q1xNd1X2SVlXilBMSCidsLeknomfh
/Rrg7a9/Cg1AXSeFAgLnd2LvXdKaOfqskYh4oJJSVd0pjJJWIgWtlPWIzlnJTdy3
KCN1rFEhCOUa1uNkBwebjijhqkJRwVtMVpv6HXVykSU82K0PLc/PknmnktYml6IT
wZIrDbaiNAWn9KVjYI1Nk/6VEdXPc3h5+kcTcvCczYO0P+1aAUn+pekgc11trjfU
pw7kU3PbyHXrTf4gb4gDzc7hYM08KTCI5lVCJyFLQdvC2F5M0tRoUMLcDYOwtizV
nVk38jQghIn4i0d1BBROtC1ITCdZDu8R12ypXM07l6LnRejWyyX6Dgsv3x0a09fG
RpX8THAN3MocM09tbRwcRDGAXqHIVFIJjKBC064tWxzI0ZLtFIcuGxSW5BU2VBzi
GMzFu1jtvURuByUGdr9UEfkV9H9b4dE3DErqmg2V1lrco+TQMwUbOgz/AOBRxwZ1
yqnDiqCdY5QvT3vc9uhomLvq3pSp0aPbxQmG+lTsI2XXcxDC8xoSMAb1G/Aqq8d4
anriud4/UoV+i7RoUF7wq+3/t6zsrwWZPq8uDflhf1DnILLu8mGI6AxZgJiHXYZ3
moz7YBXyN0y7tteyq0sFA+MoB5Efrg9sCcKQrS9kWCK+/m1bkMkv/PMw8z61285h
ppujTiZ+8vgxOp5rQ9wb+OEmEeXak/Z12+Gi753REtXJrbMRsq/TUaoSY0pxABQM
+bfyU3ov7XfYuOGM82Va1iJJqeqSOOBTK/zpROensC5RUuSxgPaP+DVuwBwIS0pW
ftvh6mVo14DXr4E+bsqlGGehiFVYetRAm/87rJgPxjcojc9dJ2Q/BflS6SObzgK4
EyjvhZh+kBYjhD+piPuKMVjqWU8sdkkrxIrxAC2oXl+aoc6HjKsXbjsrzWeUMPz0
5RJ5tPbrPa+78mgow6Wx+ofYJy+llnqtSqClCCiuZZMU1BYcEU9nUEsYmlGg1t3o
+4Q5yRmW7CiHXlkmGiFCm5S1IrrcI4K8fZ/17Pdt9PaSzIIcsQS5lXomksbLtcOw
oPGY1sv6r/OS0eio9Y9omc1VKi+LggQwMeRl2acl97DYO/RF1mEWHXmrrWlGbRLr
7XBi5+he4MIrqeBzQ8hplRXSgq97eA2qAsOCHgvEevFA/9iV0N67kdqPH25+zjEs
NfrPX3UciT8Re57CLrqKo4MI8FZRHVgx84TOpQC4ptHFzPAEUrUsSl70dN+iwaW5
7VVALp7M7+JP75MZ613JFZkIzoz2MI293dfHnh8qApDPGkE1v0GZix7vWInBNvuf
VpCH9V/9gT2qc/Gc8UsgApwZd3GHS6Om1bQd5dxv+LK4/i2h00Pjsqir32xy6etG
dnPlhiIhMCR4mf43SKLmEBP8JznCQap1NVuxNCtrQkS0SQnLCtBRfm8YS/vc2zEJ
lN1g1KwYQYNsUW9WynMPVZzFqL+eQElpIdb8sG4KWUmcI/bNHufwUK8dEN3FCxnW
/9x4EfQ78OrkU9hjT1FyRCr+hlDPOJGfvMMCkM+rqiUH0Ip8XHRV8Jsb1Z9Y0fCD
05pVAzMxQCF7WtMUot3sFqdVSmu/wckSVJ81Zn0IukUhFcXd6fo0ZpZ7Tyl/PAI0
zJMzS+uXinS84eDi11cArYKVj2G6Kraf4TLLWSmLfRSBh4gCdC2wXfPbTXSe4mBj
pt5cdErPWlyre/gD8dH1ljrj9bjkJeS12OhPTpfvvoULG99zuUv9kJ57tTFfdckE
mCzywCDBDUiEu9mTsgqD30rh2beT1mOcpywUIp5DlJFNNRGBuPAIBEku7I8jYMqc
ZYVFGBtzHAKOeYjv+9grKXrr2AHKYfXGeELDNmN6qaGS0Tt2mAxNV4dficzuh4Tm
AhGbNzS8IlCn6oVyGS80y1Sq1uaIvW+mO95Pm6vWjmL4pCa+cuIFSFVUrP5AGjBO
qf9ytBsCabE5deZo48f2PuZAl0s1XAIplyZ+BaFhvyt1VWPenNrQ0YiCeL5862uX
UcpC9ZUJTIR82Wi7MgeM26p5v1NwGYNp+N9ijeZc+gNYiPFcqXWw87Jq8LNPRSZC
UAE9u+jPGKOiAZuPigw4j8YjgBK+NyuY/eD913Kw7aINh/zBRb3oYzKfutPOMQot
QGgWhE5b54oiXNvRioB47+BCuxK94vMbCchJjn2VU3BfFvB0gqrG0OwLMD6X8Z6d
etO9d9AYBQE3yrMw46h+yujk+WgIVrbqIcfunPlLejc0+V+v15qDRRSlWcs9b7zZ
GQjlWPdVjMT8OLJRN4sJHnopzfd+GI2MQr7J95QQ3bwgjOgIkNIbSAZug5YBCDed
uu95L9KHtUh7ukyi/83npvlRTzD9tcGP+tHnf1ZEqPLMmFULtttK4Nwkzqlo9NpW
5dJyQBn5mcHvTvqU/x+KKE45+uxS+H3QiWgOOeMgJKcoUrGUhO134UGEC9pEVZK+
n+/7cHymw0Ls/bXjlv1o5d7gfCdDQ1qDb3P4E7A7ZP57FUyt7pa54f52gT/v0isF
q3xP1KQK8FxYdmFLAYaj0ZBVC8OVa4CAiFH0ucHsY/4z1rtAPMy83414yBs5NCf8
Daweb1NcVb5xQGHinyG5WEoN97A0GHK9mw64a8DS6r9yWMPj36s3zKYDwgccS+kg
QxMJiAo4A/rrUornXnbXxlORxA1tNzLa03rKLAkpPB9lsPLtwcCePXj1DDXXzFgd
6kpqWJb7JqmxukzjTDxMb0pW6ib1kGdlsjdBVCHdebdndsiRsFzut5CcylMZv8va
KG0fQYH7KiJWB1wvMzMQfwZnZFDK+jtjiD9XIt3QfXcGLHQrAWk7fNdjKau+JnP4
yioyrhskuzLfGNWeBQCvEYkA6Aq3S+Z+claI9x04gFnhFb/bRZUCEJJS3HWTEjXh
6Uhi5tWqF+T3d0CNoqY2NmGSfOtLJnDKG1MHujJZqdGrBx4Lst7GiaiF4dBOK3jr
B0iMESBhGX5OVX78L/SaVrvBN37DxD+1JXVTRQ9M79c80iSyFe4hjKni+xJtdBrK
FUjEN6Ze3QtVP8SKiFjiBeZFKyhCiuP7HMTCuD6yjSxuZUnMtlUPczqjkQgMgGGI
ESbjOg7c4IkkYIO23TMJrLMvIU/Zkv4L5DOtAEWGPb+Hi8BMR265JlJ0kal7BCqC
v2UJ1dlH078IrGOKtsjIA0vuvxp/5FeJ3F8q9zIzSw2icGmhVYnzIfuR9oLxLcyf
hVCufPPdvCNHJJnxGmc3rfqsINictpZxSUlhPMY0t/eZapWk0MazX6aXYUcBWr9T
0CKxn5JjzoBd/4YhEy4Aly/Qx5oLWkdRPwJZ4eGP5IriQCnzfeWqsrbWCV3hpO8x
J+qioud/WfUBllOvE1s6NA8diVsl4N5/j5L/E6Wp9ZRLd05u4PM74PXifnoF7v2R
FJM3q2yDjJhQneXhHAEufrCQb5lFjyGWbvk4h2z/nksy2w9zAf7+V3Njdqy8aJKa
BxB1XwzAr40sLXP1ih6rvh5eEOYnrjy9t3ZdcYuaWXdsqow1IOPrNeRIe3h5rqtv
OaWcfPsZKdkb3CPs/SkEdAwd/UI15FYtw5dz49N2qGU45cY706XZceZhEdTjso8r
CYp548yddHhwYnEzy7KWK2nsDVQrQqSh9inka03sAZLOtC4AT1wPAyXtUPUw1MD1
LS7Z747+05PUGmHxwMvqu44yKm2IxNCzN2oSNWxuRZbi2nvqMznCchi5mYMryAsF
gs8N1oIfg/v4Olhh4nkXbm/Kk4QU0mpN8Kl+9HRWqdJVVb1hxPL4J2bUmyoXHoto
xJiJV2JIC+2Qo+nHl5YNNoIgnryAjOX/EKlqp2Tc7zjDesT5BnJ+hB3QHwUq5UIP
Vonm5fd5IVHX/FbeLof40JIj3rOFRLa0wTk2KmDrZLiVPlgk/gVMVDQkSwX9Jxtw
l61itajgoKE3Qk9qLgeX+GBwYnScWshpjxsjsZ5Fwjib/hqb+ajk/tBBFvLSNzkS
Z7+IgRfb754OVeagDhtAn0LkFFUbJ8dBnQDtzg1cyZT0rw1INGc2Ub+qfBnqhGjp
rcuDMCTbFTtal264KCjxJ8oQ4f+fwAKDqz4gOR3UJPZLotdiziO4/4R0f81BCohn
vB/en+S58v6UaRLIyOL9rFSD/+xBcO8eKIPHsz9iab7iG3IuTj33gy+iuJmcQpwy
xUbDRd23H13J4z/Ae4nGv4de4NiXdyZUX5U8+yYrNdbLZNF4I9ccRI3aKbiKaLiK
1Px7mBWsxeYl4RQFznLv9q0WUld8wBcKLAQnBB3WTA56qdWyQ524MpIGFODzvi7g
VGnB4RqIczw0pcYDT1s49UrrusayIel9bLzFHExUodGX7KujtesTABceacr2WBOI
GPnKRxotSPD8Xqkqsj9QuDaEOY0dOxglxy030v+nYmXf3G/5eHq5jSLPFQqADqpM
3QrmYLyooHfRZQKHZd0FKwaP8mGEJYTsbEqF6xCAyZME9sjLi2o0FcKQfB3tjDel
X5IH6lqE+qs3gC9U+bytKdq/w7u89a3DWse3GFEWLSuADwYXFvmwFv33k70mgv5Z
Vp7q55+mv149bENRoGvh3+OSJYR7AGJmvwMOHXYZiXDpfnIAbbDD0+i91Phobu1d
g0Mkk/5maKpDbj7AbLSiDBRUESmq9MkbMGdqrUyrCAtP4zyyK0XO+4I9h+e3xdsR
/sYH2d2Tqn9wwpqzh3FVgi25JLH0VG4yjiLcQMk0NR3pRQcbj6J/xN2Jn4lxOQbD
6TwbNytEsIJ6wTiVFFtkdVz4OiOe5asQ+o1dlWGWmIks3mKLmrJas7z2NjAxK3hz
ri70Mg72RrWqG+YQFbPfGdWW2uT5BCoZvHdHUnOLSwbM9C0yRJOKfk2YIVod+tRf
iTu9OGSZrsW2WtuBrTZUvGD5JBMjBVevRgkwEc+FnHRt2Uxo7ozxAJE0YzJLeEPK
2dQ/9nTEoJuHremYRPwtH28P70SgL5ohnzayid5xHufRovkj9PxO4LNEwXr91C3U
Y9XKvPcNnxihO+QZTVtTs9kNoYLL5/KGUFMs9QZEl+QvhdW5cYOkYXJF2i59T6ws
whPqYFylUBNT0YfRnoio64tQF7NvxEvz3cw5qwrJUr3LycES/610x7qEQhCbI0vt
Ca0pLdGQFo01wmkbqDWSg5MyXsbMcMyBno8sTM9PF7PrUJ8eGbyom5Y9/HwzgZqr
AbObj0bcv0KUkJvRs6xf9q8S1W3pNx5ZJxi9wQ/A53YeOAYOtP97uKdI17WfdUjn
SXIDaKIXuNrNTqiJYHlkR63eZ9LXLjjKAa0uiJGnD8DCa0Ai4wMdEcslze1Rohb9
Uov9HhaQY5rS3h2AfivN3xasHsbU5mvyfWv64A0ijU7/EfOTzfPvwHWPKyxxuil/
eYw0JkSkQRXB/kk1mNsVNKjJ6g4MzSV0K5KMKGxbL2cWvyN6MCS5CbQosLkTr30o
5Q/ZxLfFvyG8NWMB6mh9Pbc6mAm/ivqW9Y+Yemux91OVpiLqB5Ibxc0bo7KXIz8y
WLLZxI4UYrmiU9UkvATFGf5hMaeqN0H/lzrmdUen3NWovaxSgOsI9yWrs8+dPSdl
/jO2jqP5Mh1TXYNU9yvm3ksyuJYyNJbaYMOBKH7AQgfVtydKhvl0U7lF4cc+Cb+r
Pi0jgJtaRD9jujzI4zBoY3EjFd5Iftc/TEWykMi3oRoQqMOIM5Sc5TGNndZG/t2K
EiU7GlL1SQ7bpNATGnSfcIoWNfOJm3BhOyZfLd7qryTCa25IUx4qN4dQomM18oWo
dAfY7tlSsU3s0KJXQKF73WHfrc0I4xQyWfDuHyb5QbZO34d5bSCzJA1EZpwx/Hqr
DHiAen1q7UlLxTskHQ+xdDo+FB4rvTigxqB90Bu00fh5YsfEpKkgWCDHB3HroSH0
YL/H55V12yvMnsgmaTQFmt98hL3vL8kxhCAT7Vhim9Qbbm3MQ6DKFkb33aiOheA3
spEjs//rRlcTirr3AP/mig7S/bRFWiZcnpF83P6czjxoLPRnCqpnmkA114FoGhgw
hVFAOnlY+7dJleBXSDE/hofDHhCfmfCyTei8Xvxx2ClrxWwSqpV98DH+N6f5H9ZT
kVHEZF+lFsy7lOhk3wUx97PGkhM3KiRs/M+Qu/In+O+3JEzklEI+I9tmFIoNEI0B
MY205c60lJX6QhhtOfh1UHiX0nDcdeTDkCXXIPfP7fUD2b2gfk7e5ELldVH1hcXe
k+qkS2+VjckZYZDxtm8nDDsudZtCM8RtRLcxeQHknWPyqvoWJkQNn0jGcdYMQ2d+
JNN7UF0Lb9PjMN7+hlPjP1kXote/nbjxpSuyQZ04XSsv+UQjDDZc1DdVUAqD8z0o
6s7VUhHhnDlGQPlQbDeyNSxZBEQ24XzNFuHtRUVU2M/htMz6E9p8erxoDDaO9dv/
ARDKjXJGwuCUkbglGIEmcmLpqIBH5lAIyD7HtB9o1aca9g7bEu72DYzJnmtv+eks
wzzYFPfpreXPBHWQJjVB0Aw73UODRKK7dg+aMd9o0cCPkIcoc/nQKNDaeoza5eYW
Dm9QMWD7lem91HHORUR98gZ82SjydwyuWULdpxGETNE1z9Ftz8gVBLg0bkPXP59E
S86uN9mDwZtTt0wEJv45/tHXYUE8IpvKvcFY2QvPIXT25jrJKwyoQoJHEhbaskJQ
Vn6FdQ5+H9mlztuesFv3qdzSzpy68Bu9T2rRAUdEVtsh3LSEnf2bd3+OVy9z+gxl
cgS0bw3W7KTGps5zPiJezmFt3kwS+ixzUAx+zCZcEuu4n+HxTaPh7nn/AFMte2Aw
eLgOZ8TuWyAc0gkgUNV4s27HYIbniiAD9iD48nu2krIgT2C310SNgRf15coZjqF9
WV8DJXmrKu6Vx0HD/5xSn0ujQVpPLbS53Z/GcK19Jyh8Qnl+em7CApXZFQTC/Lzl
B08+H2uvhhAKgQFGEVkQiAShKwl+6EUauvxW2m7eKSnGk+mmV5tWRAbWdIz1T9i3
LZlxGEG5e+ADGYZj9phuwBXo2GrPzCJZzfyeLyc8tlYeWzSgNubi2ZRFLgN/KVqK
i8uUMsoequMHfOBT7AwD3piwbOlIRoBA/jZC3Ko58UPOp0FbtYdpmCxodpF0UU2z
2ZDZGquZoD4lN4g51WFwC5FsIX+3vbqsAaM99a4WPIZa7io6aWcJ7Lx4kJRIE9Zu
QnTE3eztNs8x5RVZSsjnrCUEwhavRRMHGrI+6eOpDnlabFNunB5B9u/XD+eHKk3P
BRtBWvyw5RukrzgSC8ylGyPuWnNKKkwJEG7Cj0goqwby7gGDDcSvbpj8rg6nQiCz
CxT7PiJUVNvKTxcXHQs6FJhipWtMZop1MK/SB/TyqUlX5i++ZLbAOsGwAuHbdTqe
bCbRkwf6EJ81AbFaIOc2Dmu5e+c3s1C90IrFZIgVjkNc3/hd6ynsn3pbD76c6oIz
IJ2w2/98yqmVoVEzWEU9l1sTs4rkoIem/n7482amRChs3Y6+e8W0GQiiQ5WI5itH
bebuv10JSbwws0YS09ZVroAPwH31QRMx/MTcVTdxxqlMIrAyWOy18KZ1OsE3hpSx
SddmS5dqXq3S4WB+Hmoa/lbSjCJp9Jgc0sF8ElR6T1U1o9m3YeRDXZdFu8zfFq1V
MXVRiMIsGTt5rhoqbfhv7glFEoVlGwAkFKu/AjCysELbd2RODf0ZAWdUiLo2/bKb
9GsuoWEBibPbaKUxmxYdVw6C8dAMwE31eoO2cNRjBOOOsG0wpYQT+AvmMncD9CA8
XarB6aUwgrSqNPRjHzzHmlZIBcvSu3jUSkrviBZ5fNbb7YHHTQqc1wNCje2kvgyZ
qR5c3wLBDxz/Irzmku0MjayQGynFFKuANEpnsaUdB+s3NOFBfqJ7u5qOfJ70ffMQ
zmVZsxABeZU6lCbhZ3ERplCt9YTHwSlq/+mBJxbssJPybp0R0nxlYzjAZylywuAZ
DZn4Ln6zXfu2Hlj2LYFCtX5GmBrnWaVN3ufYxCuDEvb4O4pnuUyen3B4rc7+G8wa
EU7JMf/iqReY07hCVNv5qXrjActu35vBUdzbP2ojDkFE61anR4l7LjcG4zTOgG0M
bbK9rVXBpCFe6BTreMCubyqGIKVuy0YbdzqXcjHYYfXCmchLroXCsFNoGx2WWTe2
Zdq1x6kuKxhjQTrYGS8/r3IvGDcV/FPalbbrCSe+1iRKblGKxnLUwFpEU32Vr2l6
mQUpOdRKsofagFN+ktN7+Eh51M13I4Wuxbq1yYEmF2U6z40E3yN2UFNyVD8DQfaO
Mtsg16qGIsIR401mhv2Jg2PXEpxKmZe6Y8h6RJZ2HWEAcCkvA9ID6MdcttfpbMW5
fBvmqVwk443Zsh9/Hr19ze7GaL4EMgg4Z8u5FWesHBLjAPKJoqnix+xwS2ISliBs
ddv0Hpx7rn+7oxCqsH/uRNL+t5nQaoim/wkwnlCXZA6jhiwkw+KZmPs/H4MqrJdV
pTjA/N6wYPrNs4IoAlZYNTMMpBOwu+VHnji8f+X78Y+8UGK/Xy6p5K6DjYF9opx9
302cz7aISISl29ViqBhoyAoCBKt1hyrBbpWZw6PLUsuFqCLHzFEjdSQvg+BxFTWa
LIv+Oj1WT0Goka0PsLXJR69m4vYKce2GFSpP3iLmuJh4VJP8w3vR0XcSg0aZgm/T
XfTzevQ2xIR9ZQ+dfQqo18k6b0lPCUFIiNA44wR+uyvCtxtEU1hZvw5ZD0JptsYh
js3vbS8ACU8CgwRBV6JPYdPO2h+cILGqwHjPEc9JUoebu7A3TmLPwKG9Aw9Wa8Jj
UKx0LP4DFGhvdtKNv52u5+9Atf8PmqL1jrlOExEOq3il+xtzipBMYqmMUTbYSLkK
w/Gh1Ti2+ncUbFpJk5ahSClQvj68GSYUL8+yq+wCL+PPfowt3RTmNkpXT9EsyvPm
vQ0cAtOWvC4exbSJgNu+czOs8imivnBP10U+s+33isuFswpKw9hVjRRDGaWyVPPy
z1uSW3zs2DEmo/Kqf8JLOLs+2xdluoYRgIN/M6Ao/7GQNRJYSQJ+Uo9NHUWDiBdz
x/SCvaULrrp4OYymnDutVWWZVE9U3Z7va2BaG9ZxMscuKQEUGkeRaZVJfLdfCHtJ
fkM05JKTHdG8C/CnXpbo3xFCzaJeI/VL7oXqCMxwOUtLk0Zv5Xynmw91vCBz0Hqq
iFtOAyBWZBKCoxi8Ly9VNL1ciGpcEC4DvIU3HfhIrZzixT7aIKGVSWdn8+fJIpNl
tHXr2V3wQBTKTcyQlz7o0bXDSFw9qP+3poMu//PdNaiXCKi0CpQyX31yG2YWkQjZ
Gyhe4OTdIwicO5fc3AGbxWqWID3Yk4XaIdbyz9BK3Epxt5Yn4PL9rGJTIH6D2P1+
++W5A3Ly/8+9O7JnoUjgok5cC8lhAMCCVwQwF2dPtIVEzcPMTlD3f6FjJm3hkiQN
s/esAQG12Bw1BjIw9MqmxxRO8ZeyAZJWBEBVUYwQ1NmHeI4igMwkNYytXHUtGgFp
1lloYj+MMD6k2Ortf53wsHWnhIvrVIKoqWnMo+WiZkVXYYtpdRIQtM8ro2a7KnDt
GSI0ImjTSNVvBM76JPljhGS2jUA4ujGbfsJacTXHSR+Bjr7eMAs4/o1w68RfdUKF
UWBRkFx7sUKVP42uanbX6haNdB+XlkMIBUobNNWn8a1r1BDcxuyI1H8FCKNe2LFr
7jd8SDp0sTw3mMhuQi+qwHt/MZDHI0RG62uY2dmhdc8c7+RjbRlym4E+W9NMqGN2
htkdL2SGq6xsiDwnHrgf2aj+BNRJCKpo5tM8oLIf/gH19Xa6Rb1IXdkY/fpdRxCP
bt/YyLvgVr3VlQSgfjqHvbpKD/YOTr9tTu9hLoP7u82T28FRUYK2XFc7LtoOsyHr
k1Ls0SX+Ue65oM6272dNZGNxPSDgI9XDJ/OhB0MH/ijvFCbyexLd3WOC3wajPiHX
1N5B4mUAvhzNxczRpiYt5DrdoFte6IVSFx5aVHWLR4aUiTvLHyhNHEicpXhVFz7p
TtBVYu3p0Sy/jZptldjSZ0P8fmfFZd6JW1K+TuSnudK1YneeYMQJKf/b2zyCauws
OGhXh3xwQ9y/5tlMu192dPapJMUp8Wkq6cR3tI5in7XxaO4n9ZAFbqPhYOjOtXoi
2oUx789mgTwo3ktsrMRkG1+d7y21uvuEYKpYoyXokhv0j8UTe334NDtRPnAGPw13
7K+Q+p0D0s9v7ZQN97ofM5zAkAAoZg1xu06S4l+wPLPJXkQS+AJd7YYNFyFNIVNt
faHYW3sEf5p1z+f0xfqe8UZruDfRhcuI/u3NAQED2BasrB1XU/Uz9ygNpXh4rkeS
O9cL9xHNM0hb1dAMkYWZ6Yj6+2mv34gmpzvKALhbkCx4Q7UCG8ByVTlGnkBHidxh
yFqoy+rqaqgKIpuaHhC6ExbwZGW+UGK/NLnq2+/Ml7MThmf/IWdx72eMXHm0IrJ7
FnEscXr7irJ5O6v1/ZvVOagHK7cFBvPqw+x6EorcYRvHTQn1lIe3ZMp59SAMG8mx
5k65YqlBhJHyPZeyOcnNGSPJnsFM1L3ENWusRYhmg8WWovy4LT5QsGK/x47w2itZ
jSkIo8RQv8ZaDlS523r8YIQzPFqkVIVZM0DCBSjak/RGBwxs5FK8+HyEr9z8LJjc
kUlsQKUgeMBCPx4p9V6x9mQVoqpHdFU+n5h68ED1Yoa5UYmJ3/9OixHuMBgM4Grd
9WYdTVHO0yUL2hkxS2/uPCvu1H4+Dc0A3MdE29tT39hhJIL2g16rG8VhH/kY3gyT
jqlgHTfUxHHDEaX983lgLcazzjwrOIg71gSJuSyPu7sLhXhK+8kOqLDdWcmujXAn
SWRYWK6lj1rM29gcIiukfgkuc8bWDzJXwLHJgBkyjYfUVkxLmbwFrT7mN1kGVETN
3sbgq7an1MX56RF7caW0EMUTBbl9gl+DLPz73a/eUDdd8W6ctv3DGMbzWQ/UftK7
oGUM0rcDib04tGo8Kl987Rr+8vM2Ai02JVm5jBkywwUExubw2+v9AsYpCk8G2wvr
A5omGOIOuep4xOWPWevf74dS08au/V7K/l6jLQ3MeZB+bBOssdtRp1IoTDeEssVK
t6jeACIU4EMeZJ1mFOtqQmyTWDUpb3/mZr2bv8zIXzPZDIThTMlF4UMfDa2NIaoB
vOd0Dm5LX90z9ycZciOXIMEjHWUQXjfPO4jcT5L7tlBWiBJUaVeF3U88cY7TGtVN
X5lZ3NGCcX10DuuEjiOqqp4ZoENrG1eo0XNANrU5SgFKSUFZn6B5ostqwEhwAeFm
YFSN6+q8JpLxdVHnI1cNfJ9fUChOCDzfDjtwKSOrVhgymyLv3G1TBw0vC0Y+fWQy
0bnW4p6E1bsFC9TvDd6ek0vl2uU5Vm2F4q4++Qvu7A567fGkEBBgy37HmPWXqAY7
RBzV9iNJOVfWzIV3RCVZbfk267K4rMw4ax7F2QNSefQemZkWtvCo+D4LdSwtxNSW
9ZPaPSseyeMpqN8pGFkJxavcFt1lnwo4ueRtmz/hp7awPtaxvDdehj7GddtN6GVy
QoDG17BcYO3+DIL0DrzDiixuFs70qJRT+YxoNX6SzEKMnXa1c7kwt0q1NbE1zjvG
yvDob1pL33ye5TjaoK9d/DmQkERikn8JkPXW9EltMWRuW/woCbBLSCeawzb4xI0m
2wiJlo5DZveOV2pvQ5JV3N6NMuEEJ2ZyjtpiWZ+Rva25XU1aTx3pf1M37k4cvpKz
cO8JrnCwaQKpzilSKyZyae6yf2ysvfLoRod6FXtcCjvBWe65sPZV7Cj3LS5wg4Zx
bnUThSOagjDsEopCahqzbB04V3j9PiR3lLTHgqlV+TbKdzpmL5TkKtNAwpLd5CnY
3UZrDkCZUqOlH6R1j+q5ImVMK8NBMwy+h6qo7HXrM2Oa99K9P1vO+e3rXkHoD53x
LLArREu/9aXB6OnaV9Z4njeW0tMH0nYkdGuqGMvgt+Mwns9sQzsGta6iL8J/vjv/
L9eek3ShIOzPHnx/4Z6pCPkggQ/8V7ZiP6AQeL0ajdIq3MO51PxWcKc1ats9oU3G
HCGUokW6oBZOoRuhs2O4UQmZN+TCoo5VArEnMoHXMe4jW+/EJxLdIJgGItrC5jRd
TZ8Vx/mAEhmK+pXf0tr6pCbpjDyifAsdXC5W03Yqi2YUH5wjucVT2BUmYpWPpFSf
hyi1ShBbIFd8IuNa2QriKLimsZfQYkqzyDo+Ad3GQpIdnR54RXJyFRiS+xzV2Xe/
qT/UmOZ7HjwTdyf6R629Or3PJPFcCqHjwA0rIqRUSLdQJnO2MHg4lAjAvXS+uFxC
MfO9LIR5HDvI/XWtkatzOj7VX0L5y8YsX/3tAjR41st4a5plzK9VzUba4OVwW7ek
sOM81i27swjT+pcjn1cGFZ8LTstCXLVrWpX76EIlib1pg2x57sPYs/Q+YSFVvpaa
LUpdJxgiMvyHdyBtKtx8fPQzmibCw5jn7a9nmJD97PRjjNF478WxUUQ8lHJ1TJEM
2RscnkrJzgJ87WkgyIVHYbC1BcmCwIudpqClV0SNetvaBSgtfxhQnJgdd7c0ZQiY
/PfwqWmO3uKMu/hiSyEGEJnktznkCgNaEztyo28o527Ztn+vElauTFE9W8KLuMOi
HtwpasOC0p5arZA3yw9wCVOkDRvMoW0BkAxCV3bsxJKl91GAYnccDILQSv8AF4DP
6r+YFx6oKzV3z5ajfOFMA9Xg5EGLYXp4Xvxo82V2gQWWiZB65wLKY2xuLHKAEB0v
P32wHIW9eGwpzJqCsCTfJTuMcEM5gizkKvqcYTySKfq+aPu39b5b12Jp9s2CCF/4
3ZhFmpLDaOd8IPlOx2nkOpkObA8Ar5Gtt71NY6EsrM1akUUMoTjuPFUbVPSFfIM4
MOztFyzJPyIk2Exi+BxpU/l/HbqQNc2ZjRWQpfURqckG7/Us0Cd5jhlUJcVadaHu
0vMV3BtYkaFFRGcF46brFDks1zUU+tmlSstlEDyJqXYcpCKYhC3p5Ws7TF0cYcHq
VPIYY7/qhWz8hoFgPZP0953/KleDNyEyCnN5EFTNMncLOyvJDFXGjzdf8VASF/OB
WG+crDFeCSweTg3gJv6MhjS+vGu7eF4tNEDRvht0VLGnTAt5O1AHr7vgp9z+oNhC
4vI6jcE240FaUBJU7hZNpukFGtAbodDDgXBaUyzlnhByW5bpaVLMZa9EXxjzD3Ag
IJBN4pa+FieSn8MHqKX3BrqUWu3sDTNqmivn6Rm2tkLu0RomRUUrK7ns8Lk7eA00
yi2vOHn5APmTl/W4ACKLN/zQZkJIK/6BfUmN1rR6kEx0bIm2f2DyqIPtAzPCbo1Q
QfmuBApFUUXAOiRK4vQpA7nH3PsQQEGfTjotrglgRDpciaDeWqtPwRc1yd+AdbjY
QyxkS60ZE4ujrsOVVJYNNcbYqd9gkypTHpZTk0vqcCnOMObKbi87dV4gYo+uBDaq
5b5ocTMOKLt36ggfsIXGyGIG2LhUjbbnmAAIvy0SvpFC8xkqtKXwrnSOzF5IGdkp
A0qSh6GwqWMljWP/oIh9WqTSXjqawXzv/OoeQGwdqnTe2VRPAYtDsNj5hy6OG5mC
lCFjo5s8nI1iPMsv2Jcn2aNvoCoXa2cGE3ECjNjX25ElU6xW97FoiWvYcbSbh2OP
fPboHBEG7wE6YpXqGyoCf9zHmq/DFbMSDuyxE2UPA1W+AV2GEUSR4Ns6H6vbxS/r
dfPofbnDe7NxzIXr26dA3a/pnQfsgoSbRThfm3kuspcAmkt9V2G96Z3RiT9dTLwo
Ac8aQUSmM/Kt410K+F8Uc5u3c/tDbdWuAtLnSlUr7xSxg4Fm1mgYboKIMpnogjQ7
28ZMpzPdCRlznnE4C4+nNELc6HGlMF5A3at0basQkyhLQKtTq1+pJwX1lIHHmfcZ
9PM6jr/AJGbQV58kqs9pPLwdHQmdRiAvQ2lC+gD+z+Aspn5oopl65vV93jQGgSrz
EiaSBYFHPsheMKCwZRmgSMTuEE2M3ny2rC/yMzpWIaefwCIeqVWn8Xqqzl4V3JNB
MaAK1t+35zKljcwB/G0JfU0dFSQh9sZkn0vg0nNZYGXcKs9UBVpHmHkx0CDGl1GX
F3MtAmkIBqzllAhdYaCGn0+mNdW/u268ncS0xkjSSVS1t7JZTcE3qRjAqAn1IDv9
Xzoa34C9Gen4wKtfoZsOul50fKRKotTjsBawWyR2MKdZ1nVhEEi74MJlAdFxc7VH
S51VDgMQ488c4gsuzNHIAT5Peiey5O9ODX07EoaVfYzYK+gkbsrO4ATaDREHznxu
IGpowKCEAEikBgpm4jmU9PNV02nZvqROF09CbdCExEHDPV/UNlr4e7lLUHzXJT3T
4169o1ct97tWH6Jsy50ShGfZ+DDZPBz5n1JDu5Bz7IepcGTAW6t25j848hFl+P0l
o5Z1lIyP+94Qw7jPWLclzlLCj5DGXYFMZaYP5bQXDn3oK4QUoczSOrfME0wDmwaS
pDEVfVbUqLi0G8yIXGBh621BENC5OUQt/GU6HN/GFARQF6O0wL3KYuKwSFtaVZOi
doSVOXW5YxZONhwdwyRsJcNXB0ofB8V9MPTqTCDzvNyjXnYOz4XWG9nLsQ8Pcub/
OmIbFOQ2r5/AbUAGX802DUpF/8VyeJhs/QVfFTayoTuxOi0Q4dkvbO3SkS/6PMFQ
Y2P+MTTAJ6xbg2rU2j5dXT/ehNfsg4SQOaeiCfXZQCsWwZcQDQxXce2dWVoqU625
5GgQuFVAb8Lc9X1bP/SCNXyFrw7frCXuJrBx6xMzvSeSE7y2vDNYBXoXHsA6fP5g
RRmPNZK4mwtpmHWQ6DLNhTFEwncVPQW6cA5ZqJtw9eRvrsEIt2tsO1gPMNgXL3RM
cvOwQk8DwOV6csaqcsZAaMRPZWdiXWl5RQ8vilbpxFodz7wDGEcZf4B/t7DfYY5K
14KKc7sXMCQCZV1l91VZ/cRZWAM/CNSK0dWq5rr2nd5f4H9b1hf2fRc+LP4H1Yh9
1LlagLv+TsbUmrt24+AAwG0zSQeG3qWJoorhSGtQiyN3Ib769AsogW9BSHZYiQDA
E3KYCHW1emyG/mQr1l7yzKpIJrK+KcjVvJ0nuTep8LRB5Xilf0CP3WX/t0qYSSdG
N95Ggmu03b+3ZwaPAo0QagUasyrbspRqGQ4MqEoa7yEnbM+VkzUl9fehUVwGXCD8
/uE4VoyK8G2dLeJCEGcWOnMM4eZ1fHTQRUt1pJsfX1RhZYYWcrLzbSiYcbWzEywn
O21UEJyapYQRI7WLl5uYq4K1gP7LxStcS78kB58Ytx5lImiE0tkLg9+OKjkf3tWR
tgGqEEvNBaJNpbFLNs/MBI0eVGq5MvGAv//v2jtY+b8p7GW9pE77ZX78WwLwPqc9
akhZyB4fAylMge7Ps/Wxd1k/O7MjBomHbqv+NZyhaWfDozpQGwDk71KCcLbw9nRN
KYqoSFvgsQze5G69GDnoQlF8tNe6EgdqYELq9bsdG4x3UcxerSsL9EHb8NEBZYHB
Jzx4uLvAx6LewZIonSSdsZfIHi/iCysOSVF0i2Zgx0Wd6zgun3hLxrfBc4UuK341
ytywbtFwGTqieFkhs3SP27KfGDgaARnTEifb8VcCxFBiBgi2ngqcsKqHy4a2W7vh
WnJNhdO6D2f6qAhuvF0ZwwScfPgw5chisL2HW8Ze1gMYWePbleZWTd3mMlIVSXLM
w3Ch4lF+EC+JMrDrWlz9gdLNXSAREERUOWLVM6YXS8/ryHPL9BblmHvIe5gfwFsH
XDaOHsgxrU3tHuRiBuvJelb+wBaacZGVn2rIPr4GYqgcHXgDNUzXOC4IbaBwvHiF
7dMI+NsBXG1gIme4Vq0ToT4ONYfwfBSAtQDhyz56p6fzD2YKln2F50x14H7oT+LX
8LDOFbFKg/aauRc3JL0nJEBuPHYuRsxIom1FnYr88zSKK4z8a9QRhJRtxS6fXEUF
rSUe6wuRJyCGhsyDhH3nBrJEcy08fVNcPmheJoXXFnt70kv93OTxXU1Fi1Wb4YLB
r2tL8elGAcWhFutjJ2/He3dQVOrs6WaldOWb9LYHFFhoObgDIFvr7TLJshywBI91
EoC1mvH/WCePr/5ZPwPjwKVSg39T8+sEh8iQ2m5Bl2zpDU3u4WAm5RUrHkmYFYg7
XjL2ZxcjtJpsB6zhnGSxifE6OJLfWLyBd87ZUx4Pju7lu90fGCo3dfarQ3CwBVvL
338exrZChIhKE+YcgV3+VCTR4V/TDWbCoRvzeemJ3jVbUXFb7lIz1vvD2ZGr0F2h
wCytFW8fHedj/+t/Mftygr9+iO/1v/+jX2YNcNiNrf78Z1If3C0kpzAP6JZpa7qE
9k+jymLJyUv18SMxzlB0OXM3S36M+0OgO0AXLQBjd2wwUDLLYS7/g9b+bp/uvTtm
VOdnqhq3B85QD0O9yU0VVXyvpe3r8QO83LMYgxPu3ueU4LvXIt5i+jbjshXo9757
wIGYATXgipl5L2on1iCpFee52ni9Wz7MWcOPfvhzoS5VvrYJE8PArAEtc2tloOyT
38qt/AIlKNGnoXXmy646WG6dxnlDF+YV8BQ6DA7/p4eKoPzxlNwA7NMIVZ+l5y0T
LIBmD5Z1N+mwvx5nGseviftVGhCbBX5yfpYtYF1RbgvioT0+LGXTUlaZJrk9Sxht
b43g83IpJq3cyRQA37g47JZy/PpgIQtOLVDsV07bvWBJ1LkTHXAshdLk1YHpHtxF
gPzcX9vJEno8pSP+UW732VlWjeSdmFtL5p/BzexdtXE6P9kJf54xboqAMoghHdjn
0usJpaCuf/RM6558/LWc60o+S6PcxiUOCPiRmZ1YBIwgOpR2dEZAx7uViNQOIuOo
6kxuUrVr2VX2mnKRV7e6yqwFda9IYtAqfesFiS0E7uhJcDl8FtvhAIJguM9a4u3S
U+y/wICKJCEAKiQxlslKzmyr8nJ+GJjtvL137t+971Ql6xz1SLiU8bQdl9supYqc
CX0PM6OT+DK91NqYtD9kHIeEWRoZugb4J9paghIlvyeBAmMRhurlTLrJ6nDc7re4
mhQozxCMDdItcJDe0/voug57lNNrpQylvXVO05PMViQLtBVNKj6EhqcF5p1txPZB
/w+IJSkHZegbQlASeeMAbq4t51r74WePUDN/aLDMuYj1qWwBrYy+IL3/Ujgr9AY9
n3G5nL7o1154UsqAYWcD/peX/uvkTgljmT69G+MLd+GwRLq59b7TmLQizVQWeIz6
qCgjgN5FBjvzkWhQ4E/jORMN4wDVdt6c5DiC335LPhjOBT7K210c8xN8BsTDjcS/
cyWBtJyLKba0WdZO3XZSsFXDA3Iyj95NB6sRtmbh9FTeJF3BNmEcsv9lsKr4iAC6
ioURhbMS/37GPuNeNEW0K/u1pKw1P1SqL2eMBBjC4HwNpD4Hv0NjEQkiqJTvf/MD
UVIH1qD5ff93SlNQKC6XqfUl0iiefhO7rmTuKbnvxi/nWbpaVTuRYnOphKlUTh6Z
7Xm2ZBBcoYQY6YBb/VF7Y+1F9KTR7xCyqjEFzjEwBbr8nApE/nFOjWnmU1YkBVeQ
f6krxLBD3zMyM2R1PdrR0tWZ1bPpibIJ4v0i8hxJDdDyILUvytng5p66Hn7IBmlU
3YIVewHK5q2wKqnvCmJHQE5s5SJoxKWiz3ipoPz2sTTO1/wqhYZYtZur9Yt6vg0g
sgWa0Y4QkhoqSOHFo5PjcyqiEK/Dw9rDNliXhXCzOaz/8plR37B+XK2D3r3VEGMz
4HRUI291CqrpTqvAcOVJcwfwvUbqaDZtNZtQCTzexykM1o+9h06UAgizsPI3hEMD
0Z5kS+e2sKumkUNHUO0X/xXf7isjxEu0CrQidO8chaEPkqVw+6t2cdCOdTq7jmND
QhYUYn3Z1973plqlCUKbEMtXfZzRTyAKmSkbAS1rqkyYz8wAZ4ux2Kn5txHCCD8r
IxGY4i5uQSft6Ec2XK8OanonnuDOdkE56jIz+nVuHKFO1r7F4b9yXhhj8O+ZSr6b
RDLR8IwJyqq5z17ryTQbs0RpY8K7qIWPvlvYPGwhA1b/CXS+3lS0zYAzlPnPBiTI
hf6hzcAjUkYSTqWYyWgVNDoznc2viiV00sbAr4YsFH6FicWOw9qfvhRk73UDgcPk
aETVtQOHwbbRm171C6myL5nvg3tHBz0ojQGyASMGtNmkmkujjVKotTZ2cLKXmZu7
ZakVk5yfoGIZuv7HS0qSswl/gq/cvDrRULC9WIGx/96EJsr8+PcZvZHkr4UPCwLD
HsQxn9puN1zZvbGs0Em00x1u5VM5ipk2uxBDi6aGbNt6rzxgObSJ08m3EvmhoKDX
HvBDLW22lNRgAfDRtm6G5W3fRk+DdzQkG7lnFp19wLKoHwJGrfNB3yfTA5GHONeQ
8bceHdxy5GK5TijzQxqxWQMgCx/SeW7eLAD+HJmEfK/cfk5qZD8zATYPhKM1KQAG
IzkT8rdlgPnUujpK/I00yJnycjBqofWCNyylbqN29gG0nCssMmNN9batW/V/Asps
tAh2imRA0uI1bBzS0TC3ytCVQK1ai385OmdgagdpYzHe3JhXvgFXfh/+n5AD0Ev1
zi9NSybYRSIcBuRqtOKY4XjqLDWjaFwddr5eySnD2obPbhuvyMoLrKP6MpNaa0J6
wQQoy3bGy60Y0xnrqFJHDVHzaiIOzzEH8zNpCe6EVqEqlFhAnjz2UqPBttMzjovi
6V0yHr/FO421KUXo+QC4/W/TXq0gAjA9hksJF0wyqX1r0fSfAQWHVchK3HGSw1w3
opV0EYELOHkRT/qNORMxoL5DeEkqI9eDsR9dPqvMVy48hzxohE+XNqxfVcbFI+i9
iLPjLWmVFNvzwk/rLXHMmaL48K3B8Mt6Z93l3CA57qGkBPLYPFS/Z0UuGvpCsluq
fvYwnMuvYX4xrbn2Mi+z9E/bxFI5R+NpnQCFEecSdny0IZKiKfiIgIYbsrXWUTKu
3hOQP4muHga4cTzXhxmyIDJUHJG2yAFMd4cY4xlgcgvNHH5rLtrJf4fWnTYu2xQ1
OltWOo8yywh4vKffQAoboycKi0VF0TZ9TXMzU8b874JHS0azis/8mBPRpuUkY9Za
BV8WOBYLsSkFcnE8470qwqO2wPhBAJOGJEtR70xWjHbdir6FSFabd8aUPywf1a6i
mJ207JPZuuZvKHRaZuyj66YLDmfr4yCHR+IzR3LkX60NNGyh33SgnGOxZNdHN6ij
zEwaIllldEvR9q6vf+9v6l9MelxQqzESrESRHJY9APqU9xJJokV2BuyNr/JWoLAg
owkR35vP44yjCfwMqtvWopzBD9eH2FFlr1RazBsMh1JB+mcySJL+U4I3HVXHFBWc
4fLsh++PmmTJRGAtuyiDQQfyDcazsui4AOJaU7cEwfnXxuxa+ISmDV1bA2LC7otp
NzSdMw9kAiMlRuPFdb9parLLuYA8s4pziAzSbllV4rROpgWuweFtWdKXEVu91NZV
QJMeYXgl0UpcTsAX/Mqom0Vo1cg8mBj8rZiVHhhF5D10O7RSWSg1hdafo6m3am7t
KyzPPSEm1+uFnvOVXznJqNNbAbKFXSJOboDjrK9knS54TEd06xrsByv5Q2MZh4lt
6oi5k8YNmA0WwXEpn8tHf8In9Pvij+aSzlALYe6DLOyfpX0L0Fs22kbZeVmgbO7n
kte+ponQ1CLElr+qos/8iWbidQ4y8UqBONKZP31n+vRrnzTD72dMHQnZst6MgttC
pFkHakEv3miBB6XA0Ye+h3CGwHzyCfv+gVmcTiyF4xEAoFvUWDhsNZBfPbcWRo5R
j2/s5cIVuRaBvd8oQi2q9lpHzDz8OW9XRhxgOcmi0pVnigSMPZykFuKjPMrMkI1K
eAnLc2gZJS0Zu8L/7ClnQ17hk8llbVSWRA7PkX5VA7Y6k/RQfscGQz2irbVz60XK
S4iFyPmbAG7j8z0qSJGOpizV0w+xN5byRi5qapCNF78qfd5EZOpKioW7Fxa6Kfe2
9Vp6rXyxw6Q9HceI3irH3aPzRuvZmC+CDICIBF4dc4z0cYlomo9RNqVGEGBT9NNs
megqXpjRR0x4UDoSK1HnzuIjUogC6e8v8drrxk/jVCP6pTpe5dJqU9Me9fUwNRCS
IBkyxnCK7ZyYss4z7PVM5+k01FP0Au9E1OlSE/Zo53wJPhy268/bluoTHceyjdkS
Yolu7zew4LZ+T/MQAg+BNrYcDgCV4vd8Nz4f6j0bS1GWVsI4Hhn58Q9SC/oH0K6R
yetJ6buHF7ZkWwdEHuCgFe2Juzf50+VGUikz4kDcgiLCR1nFIlBZn4zV9NYd0qlU
Mz3Gl3Xn6Wm/z6EgwMg0dFwxKRrMuAQIyqs4YHOkhVhj67Z2LoRxPrjt5txln8sp
2v2JzWwb+ly62+WEUUUrtaYUUPcpiI5n3x/TkMuEIZXlyqMYHUdd7YxbrmuJRu9P
oGJanN1OZcN8RRnCVUR6fISjvWP9oge7D3q6Dy80gkseCvNollz9E1k2bqd5LgfF
NOMeieArjO5XUxTe8cbdY4sFz1bOQT+z1S93xLxhcTZCp87ZLT3jbkfNuS/rUFyi
QJcLYDkGb280QbTOHCxLTpdPPVZdGUy9NcdzdNOhNjmiL+7nGIsCPOOtcjyzkELe
rDnvK6H/lVdeWA+Qp5u4T9M/eK29eqVc/VFLG9t0/inoGw+4w6GKQ9x1sfO8+OIN
IoBXB0foWgu7f1In7gfx135DLZR5SqRxOgirzX7vA62eEzsCRNR0pl/thPwKi1Tg
+RpQerhsZ3ldiOJXcg5b7zl2rusMGOOHQ1gviqTZl+I8Ch99MuXHyxZOukwWG/z3
1gDjhWF2NxI4CpVqVqcK//PwlOXNtGlT1o00LVIlncaEAuAQHnECGra8Cfmc2JKR
Aiq+kCJH+ymmEvq7I5atwEjdbhXr9eCUMpJww2jcx4YEB9XvbUfrJVeiyRDv2Wtt
jKwIcveDgChUKswvJx56HMigOUL1YC3Ljsjr7Wve6geCST6NEkCHM+jHEtg42P4H
MYvEkdWDmFuXSQHjtdfoNgqPPwb9VuruDQqDmaadkbrtQ8pNmIMsLTsQhfoOxrM+
L2getTYpYIO7VuAz/1WjdphGJ635/EiIPeER6SoE8dD5J1KBEQk4Dryhp1NqsJVW
TAQerlBsLFZobDNBE9bPTWT/GOCHJSDqCY08gDyqF+dU9MhbPW4VzUKd2pxquh0N
kOQgrdkTsw6JB/RVNpJIZrWTLPh9MgaB7lOF7bw3cX8fLmVyO3iLmc8kB6BTEjNs
wfIBgNbaiENwYklI4n/QwgJlNvFb/OrDUu5NK8iOScmQJvjA31v3wQxsTuFREdu9
aOL89+FA7eV+THt8fHylPTggwPX+Q991yIE9+BBSStkcAEuhDmD3T2tQKqBUQOjP
rIxYpQmjPchCWVDWXDnO1QgUFjIwfPyvnb6cR6dF0woB3P8rR9qgQKewiq/ky2kA
tXGNHuCZckDQg2Ac7i2NkUrvEFdZRAJ8h3EV4TZl7zbzsFmdvXO6ogedUrr/2UZ+
D0DWJSOxOBnyV0D8wIR9HvuZx77CE0GjmTnVFHQvfTTsuV50FhjA8sL/pcPYx+25
07o2J38awGuEshQ72iQ4ObjRQp448OeB3vsUXRO4YfJbIEtaTxKpoIyMxx+M88Tu
bihae0ArRvLr76DsiadC+ONHUgs7xP9V5V1onorNU9dULUPiLLsRwj5aBWRJ3Ibu
QZDvmc16/izWei9JJvMj3GdUSmPj8bbFMm0rHrjERM6NRPHKAfWxvlYFp2xJrCtb
RM8ES8dVl0vJGX07pCQanRDoO/xqgzAlyp+dNp4s/C6kp7GcZ/dXoZacW/blorMM
71xubLY4x21HzyEruFVbWIdKzIzsQ7zK383KX5Y0KU2JXvISHlvyYsV2Y2n3QFM9
igGg8XRrBdf3oL/UMf2dWE1YPfF7m9pwFP5ltQqd25GsJcNW8DG8ITF0iaIlsWXS
QZAdpT0FpFLovKAU7ijfjMYqGQ0Pb7Ce3gzj0j8bMDGcss32LrkCI2oVJ0liqWGK
pkoGjyWY0/o/UhLMGuOz60pld/sIv9SITzGtX0/NqmCq7FCF9MI2D/XEPrM5ifM6
aSAiz/eg5F5+jeLNerRmk4eezyRRvvAeV9tkCt284yCG6psqhQwLMkQpFwALTm6I
i0OVUVUKHLU+k9rV2F8QgRmVsbfWWipLBmlp4qjtUGV9uOBJYP0XCfj4PHJFRVyG
AYrIfPNaHoHF58sV1SpTY5ntlNoHOEJ7w2IIa+9/X/34aHlZ10gnzKiPPT4zQew3
+k4nOa4Jq8C1TXYkuQhZG2ZedaQKQmDee8CgUvhi75+ZVja0Fo5/LsYnMA7NpSJJ
LrbeCPMGPe3EYBTWdjnPCXNUf0+Kcg2OqDtgKNNHNKS25KBSEA8RmzJtMr4B6EwV
9x10uGN4wf/4IfL6AeaY/+RGW3XZrE4vbPq3J7beKfSTtcA/jHI2HcQus+08MCbZ
2S4GCkZAo9hFoGBhFq3sT8hUxbxhaXwUHDSOykrjlx5KSO6pAnurNYHlFaV1S1d1
I+tha35uiVJMNuUvJ26d5UP9Ey6E6lAB7WWfAqiPZ347CIGiL+GZhWEEkKDKo2fD
rvlt2fpC9xZsNvJ4XysXef3yyP4VZTh2AJeymAGw/rOFbDckrRzVgqXLdCiGbh2R
rNoTL/2CMFzhVGuTeRA19z5hcYfouN2QDse9s+EuaPunRRr1js2qu9pTmAzQ84qz
CECVRqI2G7pdSzaYzqcmo253U+U5X3WHYmmOJa+fzfJwqqirCSHf5wRFNpPGUJIb
z3fKxspRepZOb54iFBLQhCvuPOrBmmkAkljoWB3QeCM2sFs4jI6fn0hS9Ab9NxTv
T8CrqS8brROu/S8/nIt1AEsy5Jz8SACOH0tG+mASLmFU8PH3pASP4J+z1wQojvek
/sSnfP8KcoQvyWh/5VTBEfmf4RSDGqmTfghIqdmycEjE44JELZl9fsGCRuDPkIts
C7tkkV7PUJL9eSuHOg6YBjEuKlvmqnN5qdOmB9hOmdX1N80+cIa3dklurpH970dX
mRobK+12qE7BQQL21eMkZRcuUxcOYml2YlFLcEIrH5WlYY3q9Bur5Qha4O0UJDLP
f1Z57jO3dmDSKGobucF3IilWHqROJe5cxtnUDKuiR2eahx9kGSoJakh1MNEcSNLo
ZFZ6si51J06u7yv8ay7lxKQhencKyrPYVjs992ObFYyyeb28mFjisTWby8QCMRaA
vdFaVXuK9b9eGJBo4RwCr/bhgj3RWs81sM2VAZ85M6jdEeeHdIbSU7HBSVOeAmPD
kxSThdt31ylto6QtOXqJOClXrn8BdyGaRkKs27I3v3QiHCROqphZY0Rc1lIDVI0I
E2NJpduEIJdnqFqe5DhP5vxWvZOF6OlbAH3VZySO6hTE2FXsKeNisWrBAkHM3Zyd
pHXGBufB8ZDBrRmbC9cgXkl2zKJQMT/rGDgIsXry4K15x5Lj2lx3nd2kGxXO88Jz
xlw/PXrJCX0paQxLn8NtNyTlLR0yS5hi1raIpeK7CxJkf7zCtmjd8I1g5I1OBna/
1WGcBlnuqH3dxrIXY4IcnlV9toGYlo/+108t2VUvs9Ak5PNGDkxTUnj+wBjDzilS
EY/0n3Yg34FN82JBmxeWu9RyuwlaMB3eXYbIUFYbEcYOmisinNyIfyiyf+lnNSDQ
Od/DDuuIt4Q57Si4j0IGABS6mH1shwPXAofvqdxvWqBdPVE5/k/A5VUpYjTJE+w3
8EUJhGDiAll10DNr6HxLbsGcSTd5G9iQBfAQL/Sp2INk7+tijJVURWVbhvkhORS8
CD9f7uP/i5G31bauL9mUsRlZXZs2yxvqj7OQ02TVPwSwyGcxtyra/taU5W9kRJZP
fPKW63y/8K8Iv1q9Z27aMyzKw141jIANmQtdF6JzeuHiAyMp3rt3iKph1T7yBoC4
ne+tAjv8cv10GpYN5vR/oNanUXiTmND5EomvkCYmKViBkjs7ee4iSrssRVS9uKcX
ZPEFXI14ncwNBmssDjPrkuQBYu3Zo+Z/SQT6hptuKohiLSkWKjhlbdCzOl8OqL+i
H6NpG/YFUbBAEmL1z+bS9MpYRaEnCmtC1adz05SB7nWdslNoqJ93o8P8j5w4652d
1QBRktz2sCWe8TfFR74j7wNtMKZKp8DIXGE/fVDGNHwk3xVImxUc0+5jQjFmdWLC
RFSgCmVqtS67w5cAS5fjzu5g1rak4FHSotiYHsMz3dCo1sWtl0urjtGaCSHwjIxS
gyNiaZFHfj9L7t4D+8iVkmIfyEOr4lJrab0suppO26lNAQvbP5m30wtl0TGu1ei2
aI+Ngg4AnAO9i/ahx60J2OqSkhSBuJ+sn4u9Cqq//k+ZZ8dVZ9BnvB77gYsFNEis
3egziDXdwzk78R/xjEQ4kYEuXyQ+ygVtXush4R4cGhO4m+lrZ4e1o8LmS5x/3cAV
+Iai2ZBBbnCegRxvx+Tiz/enoC8K3D43oSc7RUpYAMVKb3V2i8fBxS7Dc3NCaig9
5wptkDPNdQua1g/0CjG1nl3xjNKx5pnMQcDN7ggZo9yAVwX1zRsHcSoxRQX2qnjG
GWZj0cBgwAAzTmw18AkJrEcm2jfrClVAxOod518rl63BhspWOxopLf1Mmza712pq
ZRDXMDhhbfvR/yMFr28fruSDH9G9uyIItS64CJUaAtfDEp0BdLqt0zBFoykp6k6n
zrx/9fTAV+n9qpxfzilbUMkJXZlcAK46qIcJQgbND8oa3peVHq7h3wbFQCSlMfeU
58nVmGNSzjJ5WWNJCLqEJPizsOim5KhwXekLVHBlp9tP8uLTKOknrm63ulOl+fbX
1nDpGP+HK4XFFRDrQ1a3aa6hXtrPBwO4CTpcbkP+iyayctbEZaWzk2XJR1gYT5Av
yfQVgGAwd1k23E4MrIVBnYAN9UZHOcQLAb/N3KCpxbej4ZnZZ5MjAzSNgmwqB1g0
pd36GG28PrHbOmEd5c7Dj+RujeViZXfJb6RZYkhPc1xbvwi/y+INMJr2+oK++lsc
5JT5bNDDQo1VYs2Qdz3cIKAYhBt+oDN/DVniI8LR1+M8tLN91H2gnrL15lSDZB6c
wI2YQezIbCj56qIL4sJdJKku7+dnYXkdnwaEo+K/zWrp4iA8DJ9/psj3nmyupoJQ
wE1OiBQL79ZNZd+YERCzrLhxeZNmTkv7xJoH/UER6p3Ps1tBSeVhobN0sYiIqU3/
2yJNSjB7LHEel0px/8aRchl91jH8n3R/g+AZBWptPw0EAuQlfiSWWwAKMjh5Z/Lb
2niHrGUYr89KXhq8plpqbwDzHPzh+nAFzakssMgzIMK/jUQ1LSqXYfSZgoDYpyPo
4LnTt7FtqA/hs7HkYIF/zsXPibPeKTXmtNyy8fbIPYY7WccLa2dhqEbAr9zdbOkG
9SiSR04PK8OZwpTBKaZowDv9/lYejFNcnPJNjyQJlNIssqh+Uf894j8Zcn9mhxTf
Lv8PUDpDpl/zPt9HmKFqHIJGAXwQtlfs6DqwGXNAmuc8w+7BA1zew5FP/2Oz4o1Z
rRpuyKDHnkrX8+N3erM9F6jW/7dK+DM1stpshVf15SvDTx1GGJLLHQoKLHSYXqND
JOqARZQuBLmbBvjXZYkTly8Sb4SH1IczHqv4Y9R02mp4JdSX0fwZtQvC6NokniZt
22Ezl+JdgT15KOt2JO+Szwt6M6ZBX4V4XO21L4H/DG++eqdukM3Z9fCzPV1KF3Y2
7qQlya+VUblI9FDxeEp1aQsZhz4nA3tGGo2J4Zr0rh1Cre55gnUbOrVAUG+PvzM1
8Ix9pFAgJHOZF1sgTEKrZ/JB+ws8t7FLyGN/cKpKKqGaL/HHZ8QYaXa+kV54ERoQ
q08MVDfSDQuQ5Zy1MQaRX6CwgL8nmKnZIV3XHIvfE/eWg9RLcRB2tyU3Vs/+JfAk
S/BPGeccOmIMJXLPEwS5QAV1wNQLhvkCTvqeh1kd/JdFYGT2rTvf/pE2cwJPKSRa
W+cwZ95fcPMWtmbEDNdkyOUJSt1Kx5chyf+aRzyNLSMHncN4WxOgrDJNsAfc37Ri
m8HlNuwzVc78X2QHv8LRwFxPA/eFRtWz+/tsJBZTSerqsfJiXoh0PCZr9VpVbMgt
ns3UQssAwOIUQrKvUVOK7LJwd1JUKG3PRIj3jIMcruR1rn4Pd6H40+a4UkaZSJHF
YC7y3gv69ihHAy9haeAbopveceqZK4PnRgvMn3UlZp1S3KLENHfCemgafsES7X88
seuAwTHQTIB8bhRA38r5e266lqZ/XK8MJ3jKO5GYzKwnrIPAnkD3I8Ztj6i+PZzn
kdIs7mbd6nyY+kAHpQUtOR7FEZ8PxGGpxlmbinZIXP+7obD7G3YLVoKOYzcDVO18
ox6iKGCp/Vk3SuERgIrBvCD99u0qhlEgXyULRwQPDrxNpZD1tiKhuwANjKCzQjY+
S2AW1woiA9rRibPuDF1v0yswAaS7bhTUAKbuv1XbfzMUh1AMDHi6/mS0gQxI/xI7
IvTq9J+nayV5R4TYdkVSQZVoZ6QWFXfiMGjO3aAWR2s12Fl5Pd8Z7ZotUWpBM5uS
rjAC8P3r95Y8JBsaRjwEBeHdbXNYgBK9FaIkaqKhWGPxY+OWB3gIguMK1P+ggse9
Uwyz40JLVuX6S/zDBsyqmBlHJ9DsxsMPl9mNMlqa+r2+A+DGT3+lBPQ1P5ScoRUQ
QcVv1pH75ghpk0i0J5aLPsQ6+J1GK2IE0JUZyUERYnul7yQqiHhaJFF75jn0Qb3p
uUmkJAWUpVIoSAxxWAR7wQu8m2DxqdzHtSeeLrM4efZTGq6Y0IK4yLEDjCuuQlwa
MYE2d0ZuXMZRqQT4kYo83gnu1p+tqaCnzAWPhnTDFOf6DveF/yFuOfJ0iRC2FtvY
7+b5KWXNayeyaHq010Jpi6cInuzJWKwCmeHcpOcJAtFrK9FDz8bcKxUbLN0VgZJC
jHDcTymrDQaw1ablZad2n6Cjd3R5X/y6P2GBoR6DSVE9r3+tgJFf+3AxHeTzKcYG
t0fAqtrzQD2nWwC2P6TuHOLCoE3Hu0yPjD/NdvD+IXDZALNZ74Tb8RCIZf0e60hn
tiTno2vM4A/Kyi6P0SnkEvvJcZa85t5BLNuvbTTDSSe20dO84tiFZdTZ+rKYNS20
1nG9zwwQPOL6qqYFJwa3MWqgLwHkibQ1vr2Ya1ow/losptsRLv2ac19LScU31pIR
NQnoD++VRKX8Mne0h5QHOm5G4RqDbsWeEgFdjr6W19m7AknkzBQD7/qCWKZasDX6
JddXplbF1zcJcouTj0xDrHdyiI+DUju05zXJTtoWeGl5+N5ysaPsE5SOTJ4gavtz
JIaRB4rVHgFexobtEiI9SSLGI7boWabzlmRc+B5sOX7Iv5ThC7+fSPrZafboGlwl
BzYErhefXloQJ3lyeBVGQLOflcg+dHoaTPKs8FTg6mTC/mN9isCnBvJRkM8VwOg8
/kn6nogThbBCiBaxgfm207XfZOYJJH0OcyDwgUzy+9D4MVB8WqiOO+Q7UOIKVko6
LhCj/o0pC7xK4sU5/UEsmpFC/MAfKGz03I2VtYV6h7ZcS5sXrnrcrD9TwkTZySjB
IHN6u1lgtw+FiDkhjFUVMP4juJS/mvVIqHCqWoLnFr2VKwfAGQFReTANT/qxeYXK
0Hpb/w21LuZlzBOqQuOLdKr0EUO0BGj9mKOOTZDj9wMz4TLD9gGs22rSYA3FYqCl
agnjeRFxMh945P/HLBZe3EAP6dQc5Agy2B5kTDLZ/42bKnkbtJr+9+vrsYpNktgn
fXQfBXa4jPPH7b7wpnZwzErXunFQTdpmgBRBgSqD1gLRTlGrohFnw2D+e29HccUX
jmpELGcUBlfVX0enW9WPJMGBKUU0eDhAT8ZJPhW31jcxhujIHWxCBw7a5XmCN/pT
9jlxc5gd1blRPI0pbEA6cVjYMT2Qx13EvPQuFSTAaq5ZVpCd6lknpwsyY9jiIY6F
UKmw02ZqPQ9bOblfOi84hmg4rp261wpzEZ1A5ywc8ZE3PUUQ/30tpBJ35jBy3SWo
ndoS+k2CBps5OLJulSHjpmUANRnRLjj01bYNN0CXotim6iiI1q1GeLI1RGShwqKW
W4pBafnrAjatf8xuvhtxdFR+V6A/VX6hoD3G77BE+M6IlknDaEs2QaJHELNSXppu
2wrITtnffKANKXOutsso0TqGV4TupJuZjqGyZkwF8r62FdAZI9Dzepas+Z7ogMlR
+1LjKsqx9vKZ20Owvbqwe5mpFwCgXwyQ+FVFNYg2Lmi8CJsZhkISKbJ+oDouyOCb
Yu1+F5xIZGSKq0PGl3hDOnCLV3lY63US9soAnciMbCm7zt27z1RGQnvXaBcY9zxx
hEYPoHftr/GbAH3T8MSb/jcQ4aNzNktGlE07YpNkV6/YVVZSt/shOwhflO+UMTb1
eabiZVLocr3sfETncJHUHU3sEPtUS7iD8dZjoHWm9w2K6zzjwFMW2GBLNrq/WSTr
mNrCtCtoTsc+OImZiV3Ss2CB4ranUC7NJZOGdEUvGyycdCD8xUSgxpEYmEhgxMDr
wXDXAqIUIt0Olbe4E2Hn5RFCx9UKmY4MfeDzV0kxu6WRgqFuqyCrqq6MHwZKnZ2V
ItOEHw1BSnCJtc/uHQXE5O3EJkNQ/y/YGB8uc1aU+noe5yIkOMi0YXsNeM/8xLHn
H7hUfZBdfDM3TC2uADyJYvVJ/rl5xjaZBfOR/sTkqAVMa7/dRPxQrXo387lZyMhZ
Nics6OqHOwtqmCIJSGymZWN0mmBiOgfniyg2CeM37saJ1SSg9MmeLf/OM0sFljmT
GvaPksYl10443of6fTwiomhhnnU5giobHeCo8X8nBpeCn2goJxx3BEJomRc1+P7M
S5t4D56oJxVZHtey8UpqjAFs3/C0ifTGlsepmAebovygTcAK8mNF2mDhgo1rWpjc
Zhee9kiqM8jFmsgC0jJVVSXmTKdr5g71A4AD7cCfB3i36+o9lkinDoeSPQOTx8QX
5jicZfpnaw9KkGd9USF3X9FRRMhY5fOIM2dcK4MKROZWeeRaZ1IU3gQv+k9nDHag
CXKlZ3hdQvU77aIOlBgJgW64W734LT3Xhu3+rdcz00fUMtDmAEIKkUdK3Ct+4D+p
scBz5s7PHR0GA7UYFQVAlqJtUFRrCyOTROzBCHc6axFMAPsVjIGlgrfUhPldXgVK
9I9UThPIbyTyvvslWR9oUls0yEBCjAG0UjgoobOG9IU2DSvzkTvFlj4oZ3P4I+SC
izjRKVobuq4j1AN8BLzHjGp5tD/5B3NIpLKBNGT1SNg6LaRAmy6UI+LmL/zZcsVc
af5OImhtqGFXEleAmTv/OgFwm9rPtX1BPCyuzjkR92ZPMj5YRKKauJEdzoMKKr84
ositF//RtCJKTMEos2WJSI8tTD7+qPYdKxGZ8/Lakxnl/wT1erl1dpHXcSKErj6k
yWAeqK10eTSAPzIlzsXA37Ien/oFN+5bLCnk8rCunTfHn8eWB/1hYxb3ENBYEO8E
ZZWsOI6Ap9qDo2KkyI3ufZ84KGkXznxRphYi9tcQZUcFq6Xus3jSmgePlkJayHiF
6bKuE09EJogQsGLkVJOpe2STr8QeiONjjEzd+z9jbxAOWNFhJk6r/0Z47Qrlx6mP
GrMGunoqTzDc/6SI7QpTA14dZUZn3QKZgLA1vS1R3ZUnzOedtAZSb9PcprWhSw9b
3acB2sADyxwqU8n1mr/EcPVZsk6d+CBMKoJQE/XgDF6N8Inf0tYytsNjdXypxbz+
VTQdDjBaTMH0pVYR1GvLVviP+aG6+OOtxkbJTGwXMNEJF7kaU4C6CxAjcM1ot6gP
XiNRvZoTgjR7elL6rdUwPhgTy0zJpPfMJcqYT+tNKKISIw9vIyroVn2r06JryNXu
HwD2G506znuLHIP1ajfKIkz1E05Q1Qs2X1UWYyPwMpccG+OACZKVotpCV3LUM4Vf
TF6T8IQj/Pp9n+Tzl8+iRBchUAIVx8if8ES7yKHK6ORrDVkw6tN2NYKnPU/zyuP2
fFVNmQ+9TXlncMKYQnTVQap6YqmmPf8iktXhf+kVQqrZhkk/7u7HdcuQ0LsWJtPu
iK2XBQReS1mEkEcvGTYskbGl3KyWD+7BYCziTLEiF7uKnnGdRYrY38ZLSSTgv7cA
+mKYrGDHmtPnMs1r3FssoKjRTMxZ276Y3sDiAqxh5sIJ/GHcq/mq2AHe8Kz/u5Pj
eI2wQWABoqg6rz3qXm3EWVVQjupz0LZqfJ7M747y7y/DoELtMLh9RO+8Zaun9MMP
m70wblW0a8C28JVUXO/df0gqacqTPH3quYEBR9J9orvmSjbsC7Nktz9MEe4MzqmY
tPJFoKvQbEjJJPLQtUDzEABVBgZjFS0HY1cxVgMsHR8ej0f3n+Fy/O/R/3VqbjxP
uRpuh6p/1dJ7o181R++TKixuWpg9Hrms4Y1+p7docajMpjhHVZnWsA8ANurYeA02
+zSRZhjWYmDpoWE9KEVghbpkP5n+t0uaO8TbNOocwAaxlPKFvWOgT3hSQIHIub8O
OYsLGM571N6zW2xYBTaol8nIB8YYmFj/fQeR7ADVh3t6YP8IqLCrKFXEhoSh7H01
D38ItYpzHmzEaiDE1O66mmLe4W+dY3iRmceF93yzsSkt18P758UcdnpRTPXD9bGN
Hh8J9J1g4qzAREDC9U78XOeP6GkhBG4WrhRi2sqoYuFdNascrmbErcOuqq5zXKCS
RBIZofxDvoZQ2G7xgh7ptV+fD6RjQTXodkhwVeem2Tszqgpxy1IAau5Hhri851ZO
1YPbBJtIJczxqf42ebHyr3M4l1R6/mSukBIkKqkd18yoauDwTCw/6AVgKsFw5PS2
v4+LzQrioeVT/v8X88Do7WvpNnCCbGcj2riWkE0k0CQcquxyP0Xf0stgD0FNSEK4
KZbQigQO7TVgCkiNyXrzA1Q1OnbjNFxro+XneXKIeQrTYhLZdi/EYyqrWEpWi9xM
NlcorJL2MvobkecmglUVgsys8//nsBQAXMAaiBVFsFodkQZ6XSPSNnWGNYKmO5Ix
Brg8y7PLrt9TV+9MRbE6gb/ubkQyxic/BXenCOS+yOBWdaQaMMe/GTZxzAzBqsxX
pcVodv4kIizAupWMQ6UJd1MePN9CL2z3tOgFi/DHAwtAu/he7zzdJr4bz1/egZHb
c73q2SkMmKhBh7NMct9N/Hz3ea9CGErnjMrFQrIyPuMGaKGcoMBybc/+xc3pCKwp
4Em+5CHIAkoHfYIgp/b1R5ocn4umrWcMQEUJb2Qz71YOykgDxr0OHy9I5CrHggDK
7Txjs114hG9QL6xSA4J9orep1nqkQ1EDPd63hADhj7KYXYT67lfRe42/ZQBoVR6Z
t6mkjZI4zFe3x4FWbBhloU+y/euK8LJ25i7MpdlRuxeN5750NPMaQ/z2w1mKc/fQ
j1T7Blk9xFnAbG6c1bErSuhdE/qRH6m/8LGu1UWbCQNp1qlRRPv1rUsYUq56GPau
vEog+maHN2iJJAcaIwGsswwvM1ybnW/91uVN9CIpH7kgJbBMbsTKZItBG1Uxf93B
gVr22X3jJcvMRBw0hJvvWIcBqx5iVdkjsA00J4bqOmYffDzaBBLmAXJeBnK7Mtv5
zdWpXXdCjp9oXprIHhd6cPoakHstrdEySSllkEhEU29c1KJMLQt8xm24HWNHvrwb
RKHml5hc9/UKKcl9YuyDoILPI3JmHLgZYr+evLUnFQFg6jtW2F9JTfPdC5ruiYH4
1XR96IF6RHdS6ll1Pprvc8kqBrj+nBP+igmc3DMIXTICU8cyZD0sgWbVyJ897pK3
XkUbPhtkbNQM4hqQQTruPcFg9tKDExHf712Zqmp1ad5wVkSltlMxVMKmY7AHyQWo
18leebPhDwqEinmAqbpRcdb2QIxCFKlguNnvuF++A6VA4P3YNdaR2csIrn8sT2t5
z9n8BZEwjTIga0qQz1NqI4SAO5MmK3WLbPX3l4a/s/WqinW+aW12IG5NeAk3YXIM
ll1G/Q0PV8NofDahDZTuSNopuwdcdpDWx59fMc2x+nSK65nl5buHorR8Vtzsvo4g
ejd97gnWLevLToFVE7vp8MWQyOwHFX4K8eVtuB7YBKYpmy6etLiDrX4tic76Ns3W
KcNeFbhrO+GqUYZJ6abbZS9htn4jKv3xeglymxnC/LtdNGzXtfcNRxaO4YThP5rA
hytNps2RqeOrIDtCQcpdp7NAQBCGUgUeswiop2sk/6drqjFx2E49sVd/EbyzrUlL
wSldkjMtzL5/v07BBAbTZlZHOZ8wMHLWywrQDcIvQfuHaVdGgJNzDwQvvdgLjGxj
eLtIZYKcmDv/E4mLIx+506CDL+qZf66vCRwfijdEDj7jr8VfbD4+uxP6D5w5Z9Mi
wzzEpAiaDfc1A4p37BbC/pXseRPTLxraCpnNB3DzxMM1/28KRQ3lgglqdkqjXavl
7Ug5l5QF1gk0Gq4gdyjOKd//x/kCTr8jPiAqNrMpE13oWmpdplxJIngsU1cD5Eh7
xGLbFFju5/MGMmAhhYZaakELtDTB3mqokDp3Ynq1Yj1B1P6AJLn6TRku2YnJIjrA
7wC1P5S0ljJaooIq23l5+E6r7Qezgn1zbVyYlrRkM1QFYh5xq5BpSs/NaMokn7Rk
bLNEQZqJ402JazGLXOZ91G50rXq9SKF8Wdildevxps1aFyLx+HLxjuurHVHNYDbT
/e3L2uiHobMXqDj4Tlvd6924Otp85nVrBeFQWk/3VLfwFbv1lu4KHOXl9oBLUdQY
MiwkRGdK9/tad2tJU6oEoBfI5xu6FJk9c5A9WbSTzTVrqwdLJA0jo3KiaPyYY3bS
y2Nou7a4h1YvTavN6LzRv5EEysxvYBLVkT5BDorw6LVt9xxgGd5Qf45yxzIkqkHz
TnR/zHJ7iQ7TdrVWvaRrdBsQW8XGBm0qAPdls2+GaT4Ddlshg2GSheSjqnksTy5K
XgOjtDoTm8TZ8+Lea3/VgdtqIiUe/lXJOgo++E76pd2z0sSSe4jYqZEXXuCE9Cp4
371eb+sD/SjbYrIZJzgKSqoFM9DaiEPWPGk4LZb67zYaqLKIwROSjS1N7Sck0Bse
zQ7s8OVGJVLHym9sbT7cNVIXzM5Yzk1b5DYGdrCVOjz59hUIfHNCelrnal0h4ecl
STKvEUcX8yqSSvKTaMKhw1OTlt3dmL3dsDL9GlEezlUkjI8tt507d5DGC7J2aJmr
6IPf4XRF9qpMMoaWxhKeaaHgiLmUUzVEK/3lZg5R4DOU5Sny7mItN6vhO1BYTWQN
OQJzunPcRdCyr+y0TVxGcYi0ton3RHteIvWR6TmXz12At5c1Ikl4vXSiu1PaYEaj
ffyfnxkS11HePFP4tY3b7hhc8JbDv8LywfT1Tbc6Fy05SWCp11VD/yf5Bsk5tf4W
kjxcIjYPTp9Wws3VGQsdAiprf/w5eC++pmflx1fEAVCdjazbk6ZxlMV1KrSwxPns
F8P1EryZp8dvvruRJmM9T4OL5erAq7eNnZ3HWak7eGp80L0eoEzAi9Rl3jVQ7ahj
WacIIfYSO1WnO7JsiQL4/51dm15NiVwVz/VljIHwh6uZY87pNu+OzyirqdrNAGib
N/l6NpEc6gr/Fzeul7uxezt6rI0OrUpMmgZwgrRN4SHc3t+TySOeOuFLpIZRq7tQ
tVSKFDjEskvP7Ge48OsaQ8Kj6UiXhM8lO+X3c4qZMgajI8oMPlKJuEjIMexOIZWz
vZNigx1VEaVo8wF63RVpqNO3oDsg/7v9Nl7Oo8q1qxybeCTgfQlThdwZ1b9Oq1WP
5BgiXueE5BeaqqKYFzCfwVDHM4CPROs/LGjPf16Ag3sjyu/4h/j7i7tTa5RTVZUg
kRTY1xFoS27MACFH7qSx9rYkD+gYnTTJMF86Xnx2Bz0ZNkFcFtZU+hFM+uu5RXBY
lB9Qx2RPdJ9XGOkHGzDTrSQ8h2IlaPQLXKm548MH/QmsFHhk33g61S9oQQzMJrxD
qx8I8jRFNmhTrkwQ327Bl5M9LFPbouvqbzWbr+y818zH6ETbBcTOvtgQYZKJ9aw/
USQa/H/RKVBf1d3Of3urDsw3YP1YEe8U012RxBbwHP0+Ky5EwZLBnEa0Ugw6e2q0
OJd1NOJIF3MwW64Wz59NWiJVQJ1vsRzPEEfXpbgcXLLhxzMuxiXClgqpMCz7kvG8
xFBZk7GFgVKg+Hf1M5/BY06de3+FFgOyHnw+pQ7RExknu+XeIrvwkcH0yH+Lvkc7
AzbMgcJQwb3Vcj7/DDOJYYPFlc0T7DM81NKb4zjHN+TbTLFT2vUCdByUGslbsDMy
WBvcXak6OdCGf0CxupebaMQoP75TaB9IjBvisPe44n1exq13zfYVoWAtBHiH9RlA
s/Ac7HaxVpmfFyIxS7+oXtxksymyWi7UwYgFonBgC9uaWKY/sd2DxOLPTKeff7Q9
xO7oDlVutoE1NgPjh7fzMp79eaGhh4Noaevym6CmjM0XTHPr/U8tnyYnZXWePGnB
5TMzR7tEgzNyF0fFUWSTsNjx1QjrY8RkOVkxZMQf8yJlo+Zasee4oc7aPP81YB1g
1ODJn1yNHV7W4e9X7BjeNb6Cvx6gAiZNmGJglp4X1tNmShx07kYx9YjOr3JG1OeG
2imUwWGqDcFDXWiadbFi8JrRxpBqU/P1/MxSpX9B43P2iQRhl7pVcxSdFguyt6VG
7hyBGqjx88XiFAZYkHsrXnyp/lvAEVXyMIvngilU5nlhBVL4SWrTIpY//loar6WT
kpErD1Gw96M+KYrFDkWWrhs8SAKxl4FA4GocveJFScKT+JIZHjzOjThvvyQ/4Sga
8LYphEVGT4f17KMjd1IoGbjGJPiSddE9FQ3EWiMLLisAm0djGctnOOfKn4Y5BoLH
R6afeBpDJQdl3+x5/HBG19PeoaZgbEnI+8f04yBOseXc598ikH77JBlXmkW0uRzo
44F7PWypavbOGivRIVW0/wuZ47ztqK2drv5AQnBHPPlB3Ave4ncY0tw0T2EyT/Mr
jVbDB88zrjziCoT5ySHdxmIEcN6Drd7XBqfrZBeXgZ0wqiCujm1W2TpywoDbgebX
w04yz4GJG4py6pfc0zMlZRy4roPdvykV3uYVUD66u7FNuqoq9Fkak0qqgzHlzHd1
HfEDXFmCNQnKzJnZZdjWqCMhpXQ0YaRf9t2RxVunlL2jr++bQUr3MuO4FBuG7FpM
8zxv7L0RjWzOZ6Q8rmRKiSpL1DWJRCpNkG09w+9frUaXNDCDS0pMiBAU6ltJHQPB
vnFRKIsGSw9Be/RX0hsi3CkcRQ1VFFgNIKoIdI6o1lQqxT5K48j7X00jnB2kWJdk
vpepB5SNdFuYkDYvblUBAmQkpAUb7+Lm13zNsxF3/dsI8gzxoXbK8SHYEqeDrKsc
G2NGjeaMfzFHlei0rnR8+y1+S4tZ8cSGi7AHZpxgfuC5ZmeXzF0snDlpEtGePPi6
P11P6KDENXFVC8SSJKr3fFNYBcdCGRS4GXInvwWKJF8Dj7GrULShD6GNRAETH3tI
eKxlpf2Mdr7hiRuDJvijVxojkL+Y7hfC+p4+olZ4OETlKGHFvtLLbF/N4MUK1+Lb
MYoIAv6/QZtaf3uopN7GRSY7CbQbjDIXJ+exiPvRtHgqJgQKbmESysHbGxPx7SE0
Y5UxclGB+dR2S0aFWssFhFuv0yaJF7opWOwo+wvvb/v3r+gvHKhJHsaIVKpEqckG
O0/vZB8iUGEkhJc9chw1IzTSvU0xC/XS4ReBU3YnlI33p+jY65CM5IEB9tPHNMKU
5raLbUVXa6IwlvD+UIYDqVV6lWuLb/wthU3SGkgOgXxrua57qfYHiAJscUGrTp0h
9eemXnh+r+UFa6ZL23mGbOA4y5ojERU4B3g36dC+ItrTQ51kub9shOMeT3US7o99
CIQYFfNuIY5B/DZ64MuJCw+X6Grjlz18Fz+8v4X5NVFcu/KOd3ilD6dtTT30gXJT
iXFHiXSUVf5lwYAuluR2KW8+2vz1soBOf6FSKemriibpOIoDgReqVJmHlIIa4MvF
2cA7eRLIzLVn8S4RcNsVDtVhSsz5IfgRE1Pn1F4Pq+I8rnRout7GnWReTQMILPWe
cOeu2FGGdUZSug3FGkQsxV3VQKLYPko2kmvn2LBU5sBW8MPQW7wyKheeQsKxsDE3
KcIOZ/jlEXffKSk8wXsDTrntoT4S1Gku1p3skYet24DEUI8g1EqK/KoHi8X0wx3x
39+a/ny6akRDCvbh/p10393m+KilDYP1QLIXs4Dy6LnBYNcm+zVEvfwsVyJG1HZm
6O4bPxNYN/lo0qotCKPY4JthB3nZwZu89QArYWAqL8fg+96sPX7wQNbAOfHxq8cu
/R/PgSRqZ6COgiLleMOTSg4NF62s2UU35tLJQ82fMAliDjFdRtb+h/VONBFvjPmf
75ssF/P5934z15fzjEUKJPd9woJZZwDc+P17X7o+ddRFDaytlIrXp9UjEEW/aufe
pLX1pFmduRi2eUmNpqaoSDQMz4th37Ystuy++3KtCMCUHVWAZiwuEh8k6P/CzqZ8
mD7kobm2I3t08FySHbOr1E0oXj47efgZ9sPtS95WwBReZSSgkB8KXYBk3KqYbxfm
ANj/LIjNXXAq6rLDBtCc3+dJueDxeeKzAMwZyqQmrvA4E8oCAcx9gO3PF99WUCll
NXlu39vwRIZFBlloW2IUrReNrvL5B/AbTuRrnrFlDjqMR1hqXP0bPVE6RCf/uQLx
hqSLPEjyjmPXOezblQqd/tYRi7LyTa2jviU+0x87ivTdjX1nHrgpd/6WNfWML/QL
XyYq6prMZcSJ4lQF7k8Ae0/pqjgwxCRYyaSFeHVgzrXx8Yyd5dAjn61vn1y3XlBS
KCfxWOqnoN6w1AeobCJW9LzRMEIJRXjebTB3s92GlrXKVrcn6tuZDDXN8vQ/jAbN
+1pDsvl1zDWLaTEk4PFjFpbcDIkNfKwxSWGtGN3etpulvj2ESgkDe9WzVzEs3XKV
A1HK2z6qLItK4CNGsLjMUHERUEouOdjvn2RJnhajwVHkB92PrAgtViq2zUT4iOII
wtkuGDJ1h4au9kU1DrWH0R3o+t9Bg8U0mmf0qpkNq0Qaahqe0a0Ie53xlEcO3bGr
+xoYcXfA7Io4ow0odx+DKMxKvASOhhOIP+NsltFM1DyRCijB3ALvS35S5O6iLReZ
gnAFK5l/lrRD4pGqSab+jN2ycma/gCY2GnFdlBD9jdugKX7BLRdbfUP7J+qx1xGU
FxVtQEpxtSkeDPSt0iptcYhjE2pIkLH5aWF/uy96ZtT4zhbLjHP+kPMpHdNoMuT0
ypaZDmzhaNqyEuF4yWqcQEB/doTf4hf/YZrRT568nZb1BSIa7dtODwkQ8gbqq3YR
gN+XwmuIp9pWJlLqS7vkjbvbg8FpymCbiKiuVJS1GFt9FPIiGKNR8rpYfgU+V2zG
l+KtIyroEapaNj1rrCrmFcxWJ7iTDQGPnCoXvPQ2oMVYeWM+2fi1YeYhddIl72dY
nD7WHhlR33pTuSv5bwLUFLp493kNSVhoERgEQl5JyHCYeEOetjBOBm3sOzWXS6fI
zE+zmp/l8HTopKSNuq43VEgVvavdoe/NZNt/VN/H+8pz7/ei+HEixmvBKOxoHfn5
jlBaOaUtlN3+vLVXBF6U1ZvZSLX6j+cHcNwGLULvICEu/Q575gUnfuTdQ/NL1Fom
4GpwfpIKzjFPmOXMxilfeqFMLstzejzWy0uvf22RaLc/bESuQ9Eodu5703cdaNhh
CN9vULw3+C18fBhdAQdNfSNgYS+fUWwXWffofaBq5Z541p3hQwiDHkqzHtg8JcVZ
6hFjRcw2FV/bw5PNK8x1mQ+xxyWPEBZuNG9BdBBii1NLhMeUheix941YVlS0xtGe
bbiCRD2pBLD/FQLRb4Uva0LQKvSg5XNrcxe+cX5twhXqzDmJQZiRNsyBEbeWUKZb
DaaccPNbPNl7BPCR1kzvOnUlZ1x7OH5zI+aKxjJRhibyepbruW4vQswUy3GkLsoM
ErIL+JMxqXN9OG/Y5uTghCTS+eIaGxHEyk2lEYKXzDlHo2D5tS43mrIXXbIA8+/u
xMF1bqtTgwyBQ/TWlXVo7zfyUf4VqZMAclx5SMM11GKPFRmThntyMIZSJdBuoi5c
MlWP1LcUU5OqdGtdBNNSb1AHe+3Q3nncI710cVqX6VYIC2LFWfCJwU3Ec8dDJp6Q
8cSAnB4jeVqF/Y3cLZx3igLgzRQZR41ngo9cWcpza9ZsH4DS5ZcZ1PdSsymqHqiC
1B3iOi6ysg88uP+rgJ3BO14mPnw8G5DMBjLvOZEbDkwRiOUX1QI7HjUuMOZzFUt+
MtJCLryfWUZFMkqfki6Xraadk1aVWht+x2/UbNZAWfjAeZ8lAucljVw2aXkqxkuo
rz1VBS6lk7xuyGw5CRTEa2VacZAgmQrb8NwjS4A6Czz79frM75DXkls/Sdt9morH
I67Lolm4rRSBhnz+DPIrzxWMw4qyDDQXlVZFd4APFHFoloJIf4lB9yXZzEaX+MDu
b7+Vhso3N8FdT8V36Q5RcAybkf9WmlG+vIzr4I1Wsfb3rI/KD6hGfUG4e2ZFSNkD
Dfa5kdZNK4sOEB05aTkPIIHUS3hPwluL5XI5A7VhpmJ6KgLJNCvUq9XqUOv+mjXp
va1gsFnuVkZg0lGRjldRI5Oez5bR4JCwW/t8NXhNNkJR+gSVdhXaGhwj0LRwx/S0
xGCXfUv07+nUrHhiHwVd8WmYIGR2+0YB4HTdEM4N9YrimZISiE7Z9TBmhAOTO9uN
YraVQ07MuJF90kiTsYR2LnYTVaFbX7Xk1bG9GUIdnAmyzZwOH8I2s3jZBOnYJy4b
636dfN4y0cc7TIGrLpvhSvWHIQIgyPdCvysBbKZqLiiJSiioE5/B84k79y7SsFlf
qX1lb+w701sbEXr3kmDjfQNou1HNqVktk1mnzWCqMGNmBL9MYp/Mcx0qLV/LCIur
cBO3ocmwDX0e5q1+bX+xqLF+TGbQke8H+3r5993wjCqEGwWDh9fDEOLrC2Knz/2X
Z6dM/qFoasZTltrv7cEGzSnWELy/d7i5qNSbPlIvRqTvYDc6awCWG/pjwpkuAugZ
3ed4I42xX2Tdj3xccDov1AiUCiT1G/xdijEuIKViuKHAt7O/04KJg6I8pNMQPyfw
sChe9U4avyvPd2fPJB5c7OkQuEb/arBPOuuAkEFAVQJbbNYs29RIzRAZx7+tf4zr
3snEON96leomgMr+7NUnCxh/s3+/YQsNmLkJ6AZk9bXxBuhi3B22oGL8OZfi1V7/
JMaXCiFcKzSJmp14lhiYxwqXcpfzES+VLfn4QHFOlE8hhAZ5hOlyjln+mss4CyDo
Kn4wroq5joZWS/ZEZQtEFjT4aP2c5eQW/OmOBJMuFv+3WgzqP0qw5OrQEIBkDyvH
sV4B4EBzrgT0Rgcj4Bj8T4hN3WdQ/xC3d5OezyRn+X+pzTpMvXrcUDgiux6HoYCp
KbMNbw4BFFSCckInr+Oi5QSWJOTGXtPbd+jcE0NvZ7oumppVQ02WLUx0Jk5BQFec
v3mexMdVoXFoJKABfgqQNYfBUCkAl/dty5Qd3roH5X+NPMM5/Ayw6ygjUYUTH44T
0EqhmQ1kIuLPdp/X3s8pqd1j0SvpqDWBRLg3uZWqP3JrC3XQBE4LeGM2Uih6wjAW
xBrrwxEcIJQmJ3w7ywDjXeKgc2DzePZ4iUOABY6OmlF9lof5lZ2CkP/SjXTgcUAx
75tSDttlcu3OlEBMk5Q4wEDYcGrM0EAuTbxwIzWxaUoY0GqMl5RTJO07rAeeeIbO
V02UF/F3xgDFNhoBmKSqhm4KHA0quYnNF01KKHTv74nlkl9X3ntLEnJC/WznReko
nhwBRTKT6KwxgJz25PtcbeXaUI8OL1jgzQl/FK10mWG2nbmDx6oWpfZoj84I/nI/
kyhDk9qpW3be+Krkm6rqzO3aOjyV4m8BNOPWTmnj5OXGRB2Y4v3hxY54PN9BO3/9
eZGlUM2p062lMq3l8DX0QSTWW1+Qt10btxlwpK80A2qAzSjjGiD3tC000cK+euEF
zmuC/Z4lTkL3+31474LftPCUvbuIsVvIgT8GrgtDyVnMJNbkB7BpuQFMDvCKhe/e
s+C1fs0Yn7xqThFypNjIm1pj06jbE5JDx9y374IwNOTzkYGCr6fg5LSTPU545YPX
PVOpxJN8fp03ezJcTdHvTadWCPapzTLhlVli8Y2xRVJVejChiuEncPp0DqfQ4JzN
4/Xhn6L49O0VoeZEKg5dQlcoPs/ecEBPWVittNCtM6o2UHX1NmWllWDcyWGgsn00
vSpzOUgU5aqfZB7bghSK6LhPf+CsCIfFh+mFLogFXxqgZIPtQv3jW5A5SMncdIss
0Z00Ktvs+1wEGWt2IZplgr9njz2BIZaI9VgJunSMNgyDB/1HjZj4aAfd4hR240MC
1TQ1TO4/X/feWzWspi4GYaB9/biLt1/llJkyOs6O2U2lGEr1sLnBjUxg/Y5kBVwf
0BYzPDd2IxfoTIuRlJvdMj7hxBl2/R06Rgk+D5e6NJ1uhWGpKtngX8YTzjXkknLr
vIAgn+OsUSi16q2lqK4QFiJfWJLD+Zd6c/lvWWTc9kwbIVLpufM5ZSsB5boYISsd
VWrYL8JWUccxfQDuH1I3lUhYiNFkP/CtOvtKjXChcn/ze3hItfEufuT9YfS8X/aT
b9PYbanfOQBggBwx0bbFyEvhpepMp7dViel9Z0GkBCRRfvRFpWfh0dNrRsF51y7G
50leSz5JCL9IAxXRhSLBC40MH2zpK6t5LCe+ZyCucvHoPRf/XnBoaVwAxWYMpFcq
AcTrjdvff41UCuQgsmOKu3CYQPqsSsORBdsFAnjfz9OY/FEQReIULF421vHVkHwJ
qe/pucW/0TEklYOwtPJ9ivm6ElGHcpbWy6yrDoOEg5yztclncaboTgExzvnSs9jK
dcmuHFJSecg1+cVIXdJkxIwVYcCPllKUTgK6gg6XHInxl6j/iZb1Mz0DCJC1ZMeR
jAk0ZVcuF+7ASyZdg+zHXZdvqPOaWzTJO+e4BZ3YXrNa6hTdfGtgsQZ2T+Mu/iIz
Dw4HtkGq7xUCi8MKzAFOeXOWOjg/RNSg9ewHoBFF9s4s7smG6P1o4w7oWRVSxIp8
LxxahtXYKGeaMZ89rClu6Ho6FuzNtJjsgO+Fjd8y1WTtdNDOUXBptgO4r/YmfktW
5OO6eOR5aMt63gLwyLc/Y8o8Vj4FHFWXBmVCJLBBso8JMoyzP3ItkF0Aoq9h2naN
VihYcTaS04p7dt9blQ3mOobxoS7XZ8LrSrAzKyZcN8D7HHOi/4caw5IATXDroxFG
0JWiupgvLr10Pfu1EpzO2qEKNLxnbEkCoQbkuCOQ14R197x14OxkAywtS82jBYe7
vgvzkVaz73QC7c3zqh4wGdljdsZTDCt5hXHS+l8+1kE3YTp7plDuNTy91HX44W57
//4JlCi2UsDeet+TYTNsKnNtdM8H64nO6becL28fKtnrxWKNlXurEgyTiKOKlJhg
8r/K3xcELUrU4tHN/foMyCYGNjzQvPBkTlv3khw64z7WQ/7Vz+wlqppeDx2uXq2n
/1nbt6HCXciKQrl5VoQB2UrN1TuPYbclg92UMqdcO1fw3NulhzFdNk+dki7hMKvY
qg1AkML71PL5asBVM3w7CZf5y4e408BaJuXhib3PtUzplPSgN7dKVQULkSTs/nlz
DAlSk74RjSxN8StHFoGfUQLH+U6XsJLYGucn7jerP1+sG48jL+uegSzf/DGyXwd0
yZ79UXfmIafgGrv3PWBqEwd9Fx64ByUtVsBybSNBZeFK/Wyms/yKNQFDnx2dFh/O
jP2+g7a3LjCPgR39WZDvz3lV/80aTEKA3bnC8GlvipZ1n2Skf8rm16T0FM4a5vJw
8ITqpV3Vrvst/Ta80KfBmY58Mg9NldBguT1fyeMK9ogXstsNS03rqm2nz0q9AxXD
LBva7XYlx10UUCqlXrOh53MHzPEZzXVIrvFG6CPGGvFHvxWtjbh6Jf6MXj+G9P2V
B/qjoG3Eq2ibAJxNtlB2JYrqhRkDkQ9Qa4i0mvCRlglwVJ0AweBofmbaLqVOR4y5
bkdSEbL/peDSud7x72sVWxPT4P1f8hYtIN6eul0B9J43hCdinz3m44mcfZ8+foJm
5ZVxb4R0+pevbDa67Qv3t9dP6N956BpOcTIV3xcZuhLS/qYP+5QetkkzR7Cxoi68
t5CJBTJn3tQb7rMV3hC34Vme+8C4sMSd6+U0e4D5g3BdsNRSNq+C55tF0yO+wwUA
27mT/kZXxcjjVqei+5PjlPb83gQScyfAKP5TwhY6p268rWGFLnHNTfGywM8iMPC5
8Jwz+Q76A7NdOnQdRaluR6pVNSlqmUGjijjDQLECLmld17UzZW0dBlExgI56lOzv
+oKyDKQWyBAYDIT3Q2QodUDm5NR1/cHrSt6IJxqpQxz7cB8K5kXPcGLVoNKUym6R
dbLeuZqUmLJe+TNNA5KAi2OY/lb3IumTAeaGt0J3WTC/87km7z7hbEpWoL0HG6sz
uRk1ZSuGqFaao21HFhcNZbNsfgrqoUziGk3278e54/OJk6t3ZpkHBHpp6JL1kH4H
piuD0TpTBkU30dLP71ZvzUXVvEZeSTCL5xA9dqkqIK8kWqsQN8B89Jvy82CJ+8Za
/Zr4YJ0CZQZw97ITyOTxNJorVZ2gi5LZ8ztD6/fIQ//HgpPXHE+i1S3di+rkexmO
ab6zJbtWp3ApizLiI5k2wVkL9Ucuu3CiQi31pQpwc0F3MJWRD8p/Z/zxBBkGylmU
Z+93zIsjEPQ/Xzdhj4X5OrLNkLKi2UcjEZO0fRFSL83JFwkE6EDVZed0KMHK3y1U
rp6PvXrfl9c5h8Wfe+SHMYWCvRBPSCZQZclGaQLHH2paSTXcllrAqBIsrZbfMsCw
jsAKv7F59TOuT0guG1N/e3v56US/hEhQfOKzu4d+Nn9dlhVRD9UfugnYorxsiinA
89SQfGj4BiPyodOkrO1letLVhs+zN9GkJiKf0RC4JlKp6s83tFRvV9gzLxSBrbmS
aMGLI8Eue8RZhqqhJAChEs5T4Tkl5ODxKisJpCeLXXaCIG9n0nQ0aNF+nH5TbTNu
nDhS+tCdYAdFG/CdUsW2XHk+flDb3AbDWbU4g3AFhqN/ueAjroQxoNSREJQcuQo3
7deeBekJZqOyDQdewGCc0SMMXtQeSDVtWogJXJVramr0moMS+eYRMv4q09vnOySr
UwRGufrSA8ZjfJsbmdbOVQtGHKRD3QxlVOM5FuHVa6PVMfXvKU2TZ6gabcChkN5Y
4jwI4Fam/Ui8lBUAbc7faZUm9c71ipytl+7aLKc5892vm/SqFSFEVRsHM5F1RKd+
JiKOThH84ZxpVLK1SgeLojGTdkKPPCP6rKWLdwcj/SaGCPFXOQPrnDer1oILLIrz
AwPmYOmkRmn9+ju7HUBl7FfgZKQu3y27bhqAcNxxs0NL/fk0NyHL+cRcAh90/fr3
8HN8WnFQbGsppNWJv95joxeoMNuxfS+zkOffDsAinr6TI8Jf54Dd/a/CbUbz8LbA
E+etBezPhiNWqi1EyiQEqbgKoGlM2SUVKYAWR/UBTcDXWfcECUjFac+AFWIomRAf
nfVdVP0rG57f37IXg/gPU6Czwg+tKfTneq5WdQD/wAjk1wLvK+ZviFYeGq6Kytjc
UU/dyrVzrlinI8SEP7fCt8pn5LWpGgfcezck+WbhYrk1RYbVUEtk/nJ2j/rjjgBy
F1zejWbo9dH4b67+FGnyS3c+NzQtxCo73+Z0iYUCOh6684xDlgHjbQbIBWO56eoX
Et8YgUVytRrbTb9jMEujlm0bYhk6jIkDM2bKEcs+wqcguMAksnDDrLJY50jG2MZ3
lY78idfJ2TlXDCwSAiJURbCboYG+D37QrKPB6DlnZnNmcG3Z2TTthn3/Hr/FvrIK
ZFbSXeVYXBGYzpSOdLzlSQVIAh55IlNMOKKOqnbfoP3fogkIjNRQ27geTh8AlhIY
4uVhDxGWkWRaetU/e3NVXXyksKUXsK4SE7ubouAnAP3QjZii8uirp/+BdQ92tQqa
vdELesrEDhm+a61KxCk+zFxEqufttwCEZXOmBfC69CqD0JGOY9TSDH1TOgnZcVAQ
vYTPgc6JUtmEoJ4xTok9klfyFZggVhXArfmH6DPPHZLC1p8OUcbss5yJlntswExj
6oJT+kqYY7B1Na+1tn366KgnPAXrEb7m4de4zpjlKWk6+BKODI+OMDRqvqm/vCiK
aur8wEspEbRBylo9XTis2OdiJE06421dTCRSMdCPFZFQHkvPY2dgqLvOVhM55ou/
89aiRhyAEZf7oJCstSasR7QdPFUm8iJW4JJe0CDJeLB6Av7qJPFI05D+yIfY2B7Q
6PF3wCDY1cgiggEzCmOvam8Qx+XLSh4GebLSZIbFZtHHf6PpTHUUhXNxYzi4Dltw
PVoz39W8ksFCBQn4ecU9QLSoMvA0CaeKjeAqQCGyNrQ96nIam75sAHNSBrFRU6M8
UazvYxJVMnGerID0txcrkR6Iyq3nlqZ3LwOY5FM6ipQVxBWGPqO0Skwp012+qfvo
KNq2JaftxUSvN/vn0qDm8aIcPiJWVeUKtKkRJgy0zE2k0Ct8JcMyvKGN03wTjBvC
Hv3+PC9V3c2Jl/6WxKqaMWRiNAsinzOjyqm+5CM5i1nnUWBdhc65j8qX41IMeomF
5EtsDJnVxw8g37h4hrqf7oezGsPJOL/kXNnuPvwqvNX4PRDvNCcj+nd7gv+mJUCE
2dTp1ik0AJH9LWPOvVd37EJPE1PmquRbzqLiZUiinQ97jBn6oyh6XRFajmKoR3Kj
KzoAIU/H3BdnUDXFx1HP81C8cFRc1AaRmjhRHUbhM9SkmeY7gV9WNunVtPNwT+4t
v0ZG8aD/FusvPTxaWjBBCDEIl5ewXGTAI8O63MEh/spJtwKhfcI+K1lAjKRZWmNO
a4h2676E0Hs/+kTHS6XAyhEnxzMOWG6TsTuU4JakIYk/qtZeA1FyED2Bkbcpq73/
u4iZ61e45Q054AGyn7BvHYr57/To6ZD4viTXsWuAp7wRPCji86dGzHlLLRHwB6xK
uI41VNlIkQaZ8lprtEQmxBACDItVCLSzztrg2h6zuhjxLjSdSq++oTen6rlo0grd
9cDF7ps6r0Ru+NfXtfb6V5ozDWRho3XDNfNImVJoJqHOcP121H7UbTx9s8TsIh2C
yp8N6Kd9eM01snRow6Rf1uchDH59on+7JIN9wWLQV0UpzlgNKH6WHhJvOtJ0F0h4
+mna+gldbR+WmS8bHhfSbs0dqELAaCoyor9Q7acq+6/awpE1kAR4nxccxd0kAwle
uTsPbtNAygZ6+RKwhjoxtWe6LFbAyYDdXCINGTdi3ea4ztPwTqQt0Gxm2gR4Rd9b
IFyZZMEUTI4gK4H3Q31IbLL8BFXAsN370oxcFy/nM/t6d2tjSn4nTyUvs0W0LCG7
NgXwq/evdP5Pmb4gPmyHsxBnkJZ4HFjyMTZiXUzQxU4+KjiFDmqsOV0BHdBjRtlM
LE2Y5BBLLZTU/aRo9CYgYhDUGbsqawhTdogoWRwRlgGNX2m36Fo2q3WU+RsDs+Se
OXsmvVSb4nu6ypAbA2zoASngH+nXzDYLKUJlUDGsOoSyRI09A+q/nvBpq0xxmTdf
oGpmEcGQfk7sGXJm1g+4ISiGETWZmHXuJ+nDrc2F6n5zCzU5wBPeLzCETGWtWiDT
l1fqEcOe/ifxMI5y43UYu/IHSilkmOCIW7PACEBhLmP+NkFFJ0xCw8voWYkRJtCm
z2LujZ1/iq0PoKDwIzU549RPe6e2SJd2y/JFSxf8ofHybF9XD3gndalVQxlNWQnB
Et8xAULorvcnnHaHjQU2PH9KrFAKRMaysOrJ3pKutdZySEeTg7YQo97Im3DrATd6
NS0PSZ58kyhPgaWY3WZ7/kZ1KeYFMQJOCf4wQ2Wsq0u6A+TlPqnkDUWiE1D0p4im
/9XKaLYrjuBJqZLl2DGyyWCxXKHqaHH8vZ85YLnpFsYHa/SvD7/RJGDCEmQeDpOb
2zKtNTGZEzSqc+oEn21dqHzLa8d/gmcNuAl+H1GNeQBXPNfqSmqwDOrg+Oo5IvJF
fDtTRM2n6CfyOYzazbUCVhK2goYbobtqdoxCHZsWgC/kACmo/UVJ2tRrMfNVYAqS
ojG9CRO9Ysv3tq4fgZ5qGG74S69vWXSYycw2iinyfyMYXXMZHjTsJvw66lXT24Mj
li9+q1slwDzTfTqjsg2qrypi3LvUAhIGQXMx1i/1KuK4h1DpdtDZqI+9rKZSjnCW
/VH+lQD/1973IreuZ3a5OP6mLcm030w9v4CL2sEHbJJecacULanYNnFuQ7CJtbcn
rjKJQBShlHC2vaUa89Ii7/avvSSOCAN4xm0vLwnvHc3f+pS6y3XG4QxFfU7rTzkc
GYBIyH4y4OALdglEt7+r7g0jEVUS42Flus1lk+nuhI0d0IcpPZ4Xq2PO2Povi7Fa
s29w9FYmWC1GCG2z7WbHYL5QFIo3L9/wSU7696p7V1zk/rn/0Ht9VxkkQ3r7orJS
APQI2J2PiOEywNXYvzPnm+aLw70mm5iTOD4USIr15591RlVwCd6qBYNfCnwXBpVe
n+JHCQR9ZCkesqzXMvMkRqah4/M6ZW+kOzsFs+DwAgIk/7J6Ct21Epf2SxO9sM2D
IcSJ3Z7YLAUpXL3SE/6737y4TSdyw1LQa+QnI812jAIWFhxO5KEC4uprCOdKpP6H
VM/SpOixWlsE0Jb56FaY3XNkQ7GNbvha8mncPZ7G1JfjBu11PwLmV6RngTRS7E2n
i3cpZyAHzN52nY+HR9m0oBEpWJjmOXjlIGBK3OnXbWoLpHTrXh0g2EVwHaGCJvWV
3XoabsAtNso/GL8p+pOTjcqrHhOUzvrPIDHSnwbLcY5tbMBN+Yp94C69uQRBeMG1
7iYrj8qCCOQ9nsWZSVfP5ssVPmJ4rxo37xSo2mQRtKot8DFEKrHi/pw3uQNgqDP6
gPaIU7bms1cuTf7vkh6qRHa/xizm5P2F/gBSKxTRFx3/w7ITrMTQ4jhgcUswC06E
PIxsmyDed7LiDsEMlXm1zO+QCpPeyy5XIjbT7g0Udp6pnpj9Ur8ye05RAeIc4RIt
phqjqrGwMuaZQgRDfwe5uGQ4Aq+eMRaXQVRDZQsGAHCBaKA2utLAWSCpUefeY42B
yl9amZx9z+jedn6+pX1mSljjtYRYCXFg+in9GxiCeny09bQyu1XkJKwRPT1Im6V1
BdKCSOUHvXMFhOR+556gJNQcreHuG4Pp7tp+xGodZcYaYQcVNYbYycxi0SEyHxQ0
ouetCN++tgrRgWNbyaIOn+g0ljXfgCqdnQCQ4J0QIYZZXbyy23uSKChbGHcRs3gd
GIBCg58ElfYrAzcADrSJ4OGXi/Onx5zGHXt78cg98q/1U9nUMazSOU5sv4KrNwW1
UKVAJDwAmgURt6UcDcQ35B2nMbXqvhMRuSj/L9ILt9oEm1izkEDzluWwJ4gMyn88
3TtVMV2IiTvjh5gh9EbqAsTWpKyt5Q6TS3/OAcVSmLxN84XAz50MelzpQWWh5/GY
Hk4z/gysZWoK+z6YH2f1hS6Km0jtesDJmsNxkxbK92WuZOAUg+RQbdc3imkh7eXu
kX6eKbpGXWLUNSs9XH3XHcc3Qr5iCa21T9ONqQ0DhxKxNzWZk9bLEn4aypZgKaHA
k3/BlFnti3zLkyrFwYsoGkzPwrY6o9G/+CeXjz+1IkZG1ZIeVFyUsBpK9gdPJMTJ
gJh+QEwFCgLDXPyTDGvy1Ur/VT+nFPrYJT7pdhZg7AQV/ua45OAIOTQ58iiFlrZz
DPCmdYpBLazdONTJKIkfYdlU15KoaKy34pHEtSYbzyzpZ+RsnbBbDJfAzj2ead9T
TpFUpvwqtp7Z942VV++cl/aKkUdzga5QyVRwW0XjZqjnVdjfHcIzTNgI9Q3wSebW
L3AuxVX33pYt2E+l9HblZkj1GDSEx9dA878eBSw9GuyMkAOnEkZB79Pq31Hc+g3C
mDd1GORBU2O4VoG+oZAch9TAn5jQnrYujdKGZFpxMnKf7Va0fRdd0GywVPVSPBqo
iW22/fey2vzxGTQItMIO2J51W2JmevBDrxqNDhQaqzmW4zQXBcXtgojhmBaF2a/v
HrXrnjUljziNiiGY8nVx2r4c2oLERNnmk7q3T3zA+Vv/w8fo7m2zabGgrJgig87d
nfzBkWJ7NpBdaO9e2+m0Oq9jU4gfJK1BpGgvKZJL6VzUicYM4ZUG8v+qswzVboyy
7283aCLmj11LwJDRRnk2CMe/ibvztVkEaaagiBzosicwiWzr1KN0ywkEW74U/0fI
USgtjsQrnYr9+tkay3U4mPZTyKkeDO7h4mHJ7PA9UnA1teSv3zN5q8BUGgYId/GJ
LR8E8H/d93cm/MJLCmnBFgMCzp+rbTPiWaWz1UiCOdyhWgRwJbDmU0z546oDa11R
a3zzjKuuHuw3rbdlPZrKj3MCVyJvfRupWsNpddbiO9I4UBcIXR/CSKTacBO5pso3
EMAjT8XtG5kW3HhRSLzs+Bm9vd8y+ryd8FrxFxtX5YtQUu9JrI2d5t7mgfnprEfE
/1UXSpv0XSSvPvFQAq4z6cmNG82YJ7qCm26Jka9Aqj3T2O9yVSuqMoXgqnDl+5L8
hBPEbRYBkjhiKYVKuWnOGNVuxhJnU0njwBv6gB6iaVC8rRCSse2HDvypglxPMkBJ
ltvlY4mdLSz6QaBf/ikN2ooyxc8y1ck56uIbvgLRKfhzP0sWoSPyQBDqlUFRHDWw
/FyprNAOUud+jRAUpRlGo7IHVxKuoxgUP9ZxfazBMpTVSCIaGaMtO6BtY09TZSkv
HICOFt4mR7fm0syWNVD8dDRCzOlYm38pEgcVIbbIZgh3lT6Z6+3eawQGSCcarSeu
2qJbCQ40FJa6e8W45yT12JR+bggv3RnJAPJleUN1N27m0BQeHi735qcVo71NVfE8
wMlGiNvHGGvhl1YSr75UrT++IOb6eckNuML5kEwDiFtEB2RL6SvWjJPGOgxUJPur
i9UQQLgef+ZW4I6QO3RM48CDumwyLEA0WntGhQyYxL3ppbhksTv5DRBgXj51faPs
JLxvCHHxTSQPe5hpyun+oFS8fWUsowwXaWAxWFP1631SbqRuQJ1cea6AC5CnwKTd
UP2Hl6FIAhZgqqpnHi14asMClnTf4pIrryr3LCNtfWVIoGOA8L34X3p1eBUgUTea
UVsemANNCAO7Ij3JPiYbf3sRLPI3LTNJnOdKVyEvYdKxHUsGflc1dEI4jXrc6FnP
OT+ISf7KBhsWWZQLD9eUIvcnQe5zpAymoI2NKwN5rkooyAqOfZX8bFcV2F02yksV
03A/y7byLBGM4oe7SzClJayMVarE8oT/pFMVB7CR2da3MBqSKrdt+2xH8tyjX0+f
aCNKjsd1vfv/6/VAcQ3a69Mtl171Ubjev+afyoF+rLjyO7hVNQkTrVAvIaQjOtoi
F9OlVVOBytFr4M8qFH4QQvWTFnYADMFmYidW2THgKW1Wwmn3vVmOcPbNdnro4hny
YrN72nQDAaQOue7ZOFhRgM2YwV3MsMllelsqFPT4mjgLU52onz/ToWd/RdK3dJsM
qhf72xvMzZ0yvX7DAGYivw0mVINkMvEB23gvKt0P7JJNUPMgWuDLVLf8c9pVgQ6I
owoRmLbwCvP1P75E5jPDiChyoNW3xf2/CpbLGkqIOGmH7g2R1x/PYKhxXjSCYksh
0JyYdY0cQNnPOm3PsM1uEFTOgX+9qkplqmOaKuvpIhUMqZTvCi72DrZcyPmXfNcG
J0SZxubiehXUKrhpkPMV1LlpqCn6JmtOdb8zZfjjewTrPP1nTJAwFDpdgFMwJQws
/OOjQxU312V6cMx1tryeGRNt5vIOcAERxk0qi5JoKwuL0K3VYDBdKPlFmuJUv2t7
sHxtlRaNVycTrhMYYURVo0uIBFbsjOaXowfeWz7zwh0yM9fs2IQnIhCQ9nHtci7g
CPFz7L1x4tu5Tu0cW9QKozI8tZSNdBbI6ZA78wEX/tOA8s6F35GPcugT2KXlyIe4
oydpzSIvWbc+tH86XpsM3LCxGZpoTPCU1/SutLCvD4NZLX+PekFQR+zOOx2t+kO3
ze2UZctNV+DrdxfSdj9vIJNm/1Kesr1boOeL1NraUGM+1RqKZorWMINcTSj3lJuB
IbPwhFCSIWZQS2lIzPXyWcMMzfWBFVyUKZM4JB2QgwWMO2BM76DpbuhEqdU5ecle
IxImUNyeg6UPzim3Ndk2BhYJrtLMSBuLNEtK67NpcvtMZ4v9qO2SDWx7FPWWp08A
DtwjvYAzr/2AoYag9yokH6l2UUTwmIVDepam1/wb05jetJrjSmhVyiQir6zxuIOI
ODD4I1ytTXJ4FLtlkfYk2Iz6jE1jml22UWWpTYDXjfHrajV2aOEY8J25H2bSGoYL
J7CPfwjX6ahvf1BX6YY4vETKc1AcVAk8xaWOVH9tezXT/6MaLZ8OacOHP+EcGdZ3
yrFEFx9eXfFrccbCQ6O1I3gdunuMw88WXBKxt51mOyCNtchvUjIiQfT8t0XJAnjZ
9tJ4HDxOhgj0BJzOKS6kXZVpzIONLDL08hiTSBmAfT9L96pTjt1lriPlMqGlYk7e
LSiJhiViCKyc/W1vRTDCocoYV/KcjNCK35oxLHX+/n/gp5WR+gvw2KxMjUmshoVl
wzh54W2mFq37Ljbjf//5YmkN/T23h5psPTFLS4dJ8w2/xhdLA51JEONI/kMXABFd
pcxQ9BvMUxh9lVk4qsADVpLPxu5e49LYFxnmmrOP3GxknRTVUrDK9ZQ0QUQ7wgLu
4SpmRZsKq5EkAwaIu7lwpcXr7Smf10CZtglH+tDZ5T4wUWkyNrMpOAl0WCtatm30
zE6A9RPe+JBVRxtoFX7ppTJEajbe2xFy2k/FUdwXz3mU8SvRppfeRqeeSgq784gn
zvz1v+m242k996eSJ7vQ5EyLJszrldt3sZLpFbATSjDhGx4tUHnkOeUZhilObG7h
tp94Ayc1Oixv70QGEnHFEqBfVJpBdhRoknDmENQbx2fxbiMPtlyRxJglYKMUPVZE
cyxWwEdBZ9ZqUCQNtsxdSSen6llyc7pUbGEbWk7v2mcs6smTbA/lto/h6xS2CbA6
qnmc/zaCqhJkt9SzYyhK81YiEzPhUwzY81d76wk8tSKyuIJwqrM53UwTKYT+22FM
yJES/ZEZpdUngFCstSRpzdkA+jTPvuFJeX6eh3lKcfH6lGpN6eMgZwXjH03UAn19
iT3CPsc+MHWnD1erSNUA+1g75y3MrHoIon/FeUFZP1H63ypoBZZjF6MfK/OcIBiV
3GImy7EtQM8c0D3+82D2LiB9QNit2t6FY2Vj9Myum/5fCSTWbpljw2c63Zfw33ML
SO1Jb8XB/Rg6uX0yDBoruQ8tABo7BbuJaytNI32oK+kDIPMMN7Iw0fGILCn+OGMe
cHj4yZvmPVkf+tE6PLpedF+SeXA9QMoyXqJZpFfdkbyci15oEeDXOehRUT0fJx5k
yBqeEF0qfRLAji8qto6ObESTx5DNdE1h4LIZ0lDjxBJYhSkkMNh+WE5ie+KNl95l
VltKBf5F423GeYxiaMq/GmlqfN/fWlLC2k2wg33K7WqC6jdznKmm8X6xsVDYmL7g
1+HJp2vfbxDmRoLZxy6gJ5pnD0e1i0E5jjMXUYy7Nv10TAgH2rpQ89mhDd9SFnhV
odJlERVtkIakirImVvMMS+rhBvViuis6I9SgKUXgEcQZ+Xb8yJgkGEg08HaCFlFi
gqXhUi5uLuQaIcUEwWi98ZEpcl8GtZaO1nawEYUA5Y/vq2n3DT75D1O/N7iNRvGi
bxZvqrDt3IWk5NZ0ELxH3IYU57vLS5Fsr+jWtt2Ax+OHS7jZ+RgJFWgNqmSRX4ZT
R99D3EeMJf3QSJLX2bNI6aHk8k0bMhXj0Pv+2wqXVjcJmWEpCNG+DtSPYd2Hy7bg
HLf3STaAJikWTD9UseTVCKZ2TUYcPLoHqf9otlMHAVFoijzuV42IEq2S85iJ/fiq
NdK+A7rzfCqtkK3FT/drtpGtn6h1Qx1zb68gU7BPnFO1EwJGVjgav7ZXL93tzyAj
wmWQAWzNrIP0cX5m/LnsRhgmpszARsWEC9mKt8dI0NYPqJzsOQxu/bjfjLdvMEUu
J0vopR+5fF3AN0V1LXAD4K4/GzcFTVzv4E8W/VUzaIVnYyTVBs0lvnkpkVU65Mhi
nojybzp0mB96gslRJfj0XLEWoP0VXumYU0MbyWedEyeO0orW55XktWiQr+gjLSSs
UrOq9U9Hk2PNnEI7fOKXUcaoge9eIk+JfmvZ0dl4J9K36sP1DlaP4CejlRTE34Sg
h+yCedrck/4MJyVXbsprq9TcCmwfTq3YlJQWFHDswmdDkHx9yzpol3HZLNwpwYkP
mWR/C8QdiN+eo7JY71nqsx2OfJAUGW4JT6kxWETNdjhTl/xXhyon6SqQpwHEeFV4
/06XokIb/0rQeu6YGSdgAGne3a5RjCw/XCW6iSKlLkpkChpucfMHKgKhDe+H1zFx
ATwNv0nD/E7zCdNiA9jtxEL7E+s5UHbQ08ZrqvED6HmxBcNn2VXvJVDdU3jz+/74
/Y9sFNbirSxIdbscny+plYHtnydfMq56pb8R3D60J4uwkYN+r0vVM8J2fPqrMAMe
HaXf55i913GxQUJxV3IWCfmvSyfm0aeHZ6aYAdkyIIMKz5j/6ls/mpClZvsdccT+
VM9fmsV79UBIiF9EUdAdUV9SYf2oXCrVBL2aqc1voi1b0LZF3t1bQWu+oNm9LZbw
UkwMgXXPDWxPlpGR0jWCpHuEDaemLEDfzOuQCe4MWAGBJm0T402+KDCY9jNMVCEM
gmJQeWevhfOOH1VQZBcmGZ68cxT9CfOAMtZ/60M0BplKtc5n9eVr7MmOG/X1zcO0
5rHTiFdoODbOGKyZ5fpCflOrPvuGMX6raDPqpVRx1E47q+gjZWpT+6F22WVlg7TY
JCYiK/L4O7KDaXK0E8wv67UscP7tW9zgyO9FoLUpFuvf0SIKo/z0Lc6q1rhISX69
VmnLC9/oZISlWubG63StwRypsk2tLMJQYOl30DlUOIKMUYzcu2vpvBCfGwQsMzGJ
cSfGhNk865DdmIxQKa4lG6J7/lSk16jfwo7QRh4yMvzilfySad8mtAmuvcobtNaC
HF00ZdR4ElqqvN3BxDnU6TTe+0XMmEX62Jc5nnuEzX30SwAGzirUgc13aYE8lUBR
zFpIp+fJoG57c3hV46CsLYnxF5VnMTRey6/bKdHBfjGSTmsZUBUZtWtzTxE7fKPW
XZ1Lhicdqu6qPhhdwrgw4NfFEPDXj+BbhdXVKag2C1KUGYzJq4u+lpuEa1m7WLKi
WMWWbesMZf+Aaz2Du5tQre0qSSIkQbC8eqh/jZA3QeFpMtJpr9c5D4HT+3fO8JgL
k3q5u65sZFaz5rpGNgSU9Q99EvDVdEfiID2enT2lG8LSDiVnL/NayD6sx0KE1lQl
ZheAdGVL2/bHR2H7g6rGf5CxzwNdMdQLFNWJG+Dly0/ovnOLLC6GAGrpAXa1VD9c
zCRQjPCpaKGfBMSIkdMF7Hg0PUZ75ClPwqKIuMzD0uOl/X47s5mELzTaQ/08gEpp
cs4XEhW2fy+k+6eBS7YkIBqWUcIHRZFA+aDN3zO0wRWNt5qlFk6Cei/TNzI2I8Wd
EY2h+3TA9aOHCci24lpaBDHGGMVYJDsjaPG68W0kLNORsAqLQOB5mRWkghpjiOoS
s7xEmBglICaHGXwxyCT3y/DWKwXtXqCora2DkD9DI9FtNrZ2+4RlPPlyhZOjyaRY
gV96cV7eD5nLE2rF4jpBfIghQ7jfOytJJ0WLUsMtuKHmm6AStauChsxEm2fmahBj
zq4nr9mE8TBXocqXkU/S8kGIvMO5NE4mDdlcaDGsx89MYmM0tL4/uQ6crA0TR1Hf
O2tSV2Ffc3fmjw0zQSA+sVk0H1Q72MP9Z0B1AD0a/O/N4gVy+ikhqc2P7Eoi7www
hxiRog/vi6CY6VvBsCvKij5YmwCED0c+uH7UQ1zPSPNDpBKQGqrUu62nSdycz6Qa
mOPtrmUhIL+RJrfWeGB2eqoqqvmGT1+v2KiQAepbqm1WDHHl3dWHIsDt9aq0Dwjd
51GOmChROUZhCM7SndeRCwn2j8s5f1bL4CHOuJE5gKynlmvXCcxFVRgFNXoJ7cV2
28xoThB4WgriQqVpsRFkn1bsCE6JtcHJCAGEU4hmgAfZbcBGpP+K3bbjswGoOokc
2cxmRLHhPp864YIhyk5GdpRaT8lG43UNcCpFwSlf+SXktBqiBaoK0UiyW6ChT+H7
2Y6gYj5zn+ZeWXPr8V3Gx5awalQgeWpsv+H4euWIXpRzqvl3jMNPXk98SoKcyvUP
MtzYy+z/WJasctpsHk00u3OvZA0WD2Jv8lt54WzqhccIFKtSdMau5ql78yVp0MXT
v+eN31WcmUgjWTsbUCjaoqvuAi7RKNdCisSf6UarsfzL2nb+7+R/WzetfKw2HDca
GqVn13dRnbm7u4vCwFnXpF/0s1XKM0KPodXZVJ3VKnMWgWq4sa5p+kQhsHXIr9ko
6ALVbgTKYweDRkjOXGPITN65Mpgd08YYtfdjNuJ66qL0su0r/jhpy8QRCFtr99Mg
DjDm3nGgJ4MjtLPQ+Ak/RfDElu+KNRPP9OuU+RibCZixN1PK96X3d8jS4q40gLNb
k3dEg1oaMblPzj5HNYsGxMSvszvaLpLHX6WVp4gV+HW9JXZT4ZYIKVeHWRcXidS2
Duy9YR1yF+QApwZ5cmTNymQPz8aDqRFiEwvwswVq623G7waY6t1/I/z/51YB7BNW
HFr7qiksDBWIuNxqiatkSIUTOCekhnih7iotHHCh5ZG4kPNoMKoJzmMFHTSDuSgL
92EPLG4dLJxzsFtATXUMG10tabRkG1ZLmibpwQSleXiRKVNSv5DHojECykgqLaz6
deCX3LqLANRE/PnynwBAunEngmcVZo/UkSnP9k3D/64DBAKB8T/LmRXiBM3f9Jbb
meGS69yjaNysoAoLYRLD7A8sshXRUS+6rongZvWXel3TYmU2bUUj8oJK6pXvL644
V//IX6l0gJG3esuHkBu/qHvF6eaCaFs0YHKfVgUv7dtc+izSbe2Xl9sMs8nCppOX
52Gdwvs0JKOBPZ6DI38FJpXy8vBFbM1Xk6Rlk9yXvF5mDRHKcOGm5FbrNv8ZR5mo
HnhYYvZomWSbfc07l58aln+yh47su5/wfRPekhCbq5rZKCuRZpC6YCRi8Wvpt788
CnwtqUIaqR7k1VihRcqxbTvKqwpnL6zK6D+sGfzPS/V+fG0z3hX3sWV+ClcXyGjV
HieKSBfmmI4PQBA3mtqXZ3KX8lFPyX+wULRnIx52QntC5U0SnihNX+GavarMltLv
BO+EoRmHKJI0OcEjU0R/6l0ON7X+K8SvsrzR2m7DlTj3WPBTvMB5VDv5eVbc8Wqn
wBsFfxS8hQnnaHHhFhdthlplQ0AAn4mD1vUi2sqLcbfyqp1ZXdRHa7yJYdy3A9l5
pNzGu4JTnAcvw9CtPVI2K4aCOZp1OwDOW2YufNXKrWWT+CgjhGa14xsuOftrLZoy
ZLSdhaTQNScsX1qhLo6nGUBPr2f3U4RtxSacv9xMdb4pi+LskLTeBC9dhBRhh5+n
7r3Zxj1Xwar675xpRpg8Ne6JpgQ35JepvN14uJ0tixBmfUlwp2BPUDnKtiC15hHu
QSVaC+BGq8aEwPkVUt5iEmEHKpV37QMdrt94GsSiDy5Eimj8MRTf4ACVzGnLwHPE
c5r0mszBafT0asHg9uTGNgZKQ3jT0lgWO6EBKmp8SSxMJqwq9N0e53fCwn/cTJYT
zZ/XzIsaXQIduMUGCmAzd1nN9EinGmXEVe/QbFXXmfav/MI+DPJHIbfBm7MK7gy/
v0XtLVFoS/yiwiPhKe09D59tsO4b4gWULwBwX9YC/PLPHZXxQVvSUa2oBPJTPvDV
wHIqFfUjbIg1gVNSnRUag4kf0+BIV/jAnKrHvecmxFFf8Iz/Y0bVAExylIMhAFnY
nctZPF4HE6OD3+Oi0NZC8iKu2kA4cjeHeBFST+2mQW1aW0yEVAwZtJsp52VqpEVq
U66UrAdC3CGb02br19dPQwaktbeBeGLtjeKyMyoA/+nq1Op1PbannvBrAX9PqJRZ
wAzEoM38wRMaf3u805BGD8gDKttUmIOU+poGPtSXn2kVOu3ieBLO6u3dztKe9mGY
F5X0Zejb2b/Vh/j8rFMZN1+KltkGPp46gdABn/Y9YUWsrKiyBiGWk6PaRghhYQfb
GHOBSSp1f9g/Dlpla8CaOkeJ34c4EW2ro8LFzn70nB9WXIVyPDQMPC1D4sbDQEC5
zqt99GmH00ZsmKLifueA+VtadUr9ppu0YqyhTUGBcOPusb70PWwiqNBWmeTj0thU
btkPFXta459mu8vmCMYXDVoj7S15TXJ3B70lkn/+wmH4lvqSLz3Lu5+U/uxvS8Et
0g1KMsLu786eRd4zkiOZgjNz/WNDHMBcYD/3MphB4hhd9cyHpM9OyH1MvdEV+h3z
oS57CLoBxhaFeZqw1IPY7pyeVPzPGTEDqyf7SQ4y53vcvc/tnU+HprcedVNtEaP0
B/qDSU9s56G5fE3iVbCI8gSjJajhLFCwSdHB/amyDOUoFEH4GNq9zFKJ0sjiANvT
feEauZiGrPBRIpoZ6AZ5/o1AUAcaPx6KBW0gQazIWwyNvpKV80UVe+o0gd2xJ7tc
e0aAE7WgtGaSRYCJV4UDu1rGI6+tjNskPe9HVU3C0SeQnDz5OGPZm7TocgF/NUrh
zzhVSj5WoroP7a+J5thJV0UHrN7076Yfvt8doCEbvH9oWOwU1A6D3dqkC3BwfPWc
I9geyumtf4e+TkYadG6fu7DPydW0uWg0ETvPyNJkAxfiC0orV/LognoOb8Msf35O
riMSAPGvSIFX2zM/KCQNN3F5M20fhqL+IkBOoaBUkyO4nGKYWzELG8g0XgVqW+QE
K2lLocdc0WnsAenhwno+WYAiLc5NgmZKVrahpMpegdA79ZmzKVTr95QPaXuGb+ic
KmY9JYj8zsZ9zpJhtCEfcs6+dt8vtqIFNQ/bPub4r8VmoftpsWQgsiOvmtRPQoX1
GUfJHcgzekexuLCdm0SNTde5DhDhMu1O3AZKpSNm8vNFtH7FNhIyxm+xkdAzJHaz
eQmqFAszKgtb6kjO23DUPgZt4hzSD0LsnKeMQAjjno90WoYgpcdJwkWDkhTmtYC0
RgCvTZ1U8WI4WOr2mrghsJ5yCVG0Ow5lsIUEuWb6EU/BWClGuwPz1CZqwoUuqij3
/aDA4P7T+v+zlk0+hQOQO+ynYPkl+xxo+w3Uzi06zsify5U3ByoixqEJPfij+HQ5
kWR0vSaGc+n2mvUqtNVS3/yu6Tlbc+1w/sDj1QLVV5/5fLi1I5Czcup0B2EMA3P4
toc1jD/L3dJbUdeuZ7Qw4sjdqrZpgnvN3WPPXqXMnRST54CNfc49bjO+vQkrkoPK
NyCG5ZqGhTusonopznquXsE6E3hpDtpFGoc5jhswx0OrqU5shRRVDT08AcDMgRwp
8NsMbAYXXABr3sOQxXRnYitPVEa5D1dbXWoyri3/vHiYP4z2ZZg2UKwkxQGwxmGu
q5n1zTS1vkSk3CGj0wpRHnU5wML+j7KHOXSm0nub6O1S0Es9HlkzJor+rRxOuTym
xYIQ9B5R/WMAHuE7UN8VzEsSnHplS9Hdk46cyncfXam0ARgNzki/6QZrZHJXoINL
AGiqHDUFF2arEY/moIaX9O5YzaoGF0NFXmZi8tiW39hwi3XBERX1vEorOSzHxHd1
U1NliomylbJ3+msq5cPOFc4c5J/xPJBfxxYbngrs3pMreFrMvvQoRCUfrrda5QTD
Bzh9LqA1Vq1ewYg+fhUijci8+Bx8ye9TDJTIKDlHEq0d1YbGX4Mpb9UCMZXcKLFN
0wtvEF0fYQpuiXrroFU3k9CwuyuBATsBmWl8UaxAxA4UqmDzeNL2wfHMW+8LDHHb
ct/e3+zCFoVQj8c4wVj7+GLEptg+Uby8JKqeq4hpJ5KiKMtChkHZuZPRFJ7g0qcd
JLCMe3Nz6hEMadBVuPjmdm/hGcDygmGf2QKIHZ1YYvtZZrucvys8kaDiYsq5vxcF
RhDT0Qck7n7o2UZNXpmLAUkwFHUU7PvtKYhBO0fBbmYxHYQSBsg+0us9IFKRjYPO
gTiKaCHBsqnlLvxSi+NBWzs1uOOd7DsEmLXfCe7LWFpAY6NSdtTDEOAW5EiT57aC
qUhih+vKkVxSy75Hy1p3GlE56haBLRNzahOc2MxAusurGriGatWq0iH2MmsBi/GI
pktFn37NcmNpFAvOp41kVdTVrRNCkC40H1tq46bPUhDvW1e4mVglja07kjMB5IPm
x6FReSUEX+6HPYZnXdCnDbUfTjMGr+A0f5c8ayr6g88chVte4DBs9a+YAloMWVgr
STkCSTtBdev3ZxHpB7Rk+c4fukA6J6IIHMqn/twkqm+pg6kzos5xGXgYAfgxkjEb
X5ovoJdl2QcbFDkwrBVtJAJ178RNg5CcQK6u7Xp4iqhdN+7EUfm/CbcSV32dm6wu
wfmfKkdwkFX2JSV74wn295PclK78h9DNMCzSig5OZAuU0xEvtVspXiqd/DUSQcvu
kNKOM00vb39wp9EvDQaP5aTflX9WvS3LhCm7q05rY+m+oSCw5+6plYlSebiw2KlC
8KG7DYAvUJweT4CUAkshh1pgJk2RDEst1dCqk+3/5M+3Pn2tI/yj2GeurkFjmTp8
StmXJlaUffAnpupmPl8plYKN+W/87h/vBMuh1qRvwd5AEKHI516vobm9fgIOzgFw
elo1EQecXU3FFTcQ4CIdlnpvf9cANP42Z6edq0wgxB81JfaSLyaXTEyVvOOxAXYT
maW1ju9g9+DDALloyejWdL1yQ5JeufxgB324MjrT5VHpIqX8IbWTeOAyGmRufKcA
OSg3XdTo93A+BN1dZXhFT5xK0wrbINkl1yVBBxBqVZ7ywjOWYl2wF1WEKH37RO8K
YEuTKRZGlTq0wncyzHFpjs36l/jX1aVTvkcHPs0gErfKYr1se0pxb8sDUg/8J4ln
stWSwYPTHVhlvPBpXTVbihnf7byfQibbnnh9Y2d9A6LEaODbctj05MPN3VnVBxTd
/i3TLw7X/QyseUT2wQhB7dMn8nx0dcDSq5kCeRyi6800ym35hKCPf9JUxPCAd+UZ
fOEkilpZI39ZFryqlFHnbWvy+rPN1EgZuWBpJ/p2Sg39HhiG5pAR4669MOFZZQiZ
zWUMLmVRlB9st93Rqkwn2QtH1z4bfp6D2uEP93ZkosKHerQWMwC+DD9GqDlCtZMQ
foMQ5iUoRFxQQX0X25/6v7ACLQgpB0xfruAE1mHY3lNmfoB3nVhNsWMq1GcvMCtS
sKK1EbRjJRIrMmgAlJXEZLNYuNaEyabc7oAjIVx9Rk538O6pBQx4ItV30WyAOBy9
HSl9K3kSAP4pzlzsR3AoL7B+DTgKoUdJaa6Swn8whvoHpvCMUlI2YQw/nmbjd20u
QK2p/1wm+9kJaYQrCGvzut5kNFMYErjsrnh6gZSovvW/ift0hjLR/JPyDcxAuqqW
XK4sHvJFDMvQvmxg4uRBaRSbm+Br0I0uYEwQZeJnkUUR6fesdr9h2q6OzF2lnjoG
N1PBpwWA+K8yR5r55mPvSg4Ayj5H0PdCtiCosgEALSNy9uScbdl3sm7CUJC54D4K
xitTHzeLBKM4WpDJ3LrSQHrJ8FNYqQu2IRRgUjOyNxMLItcpN0/Ce2N/Gzmpgwep
PhRhhM4qOD4TGacDr12w6RyVnhkhEO5/BFJ+k4trQc4j0rXPx8s0j6PDI1xxhCQS
cPRtIRvXA9vcWXK5CK+NneV4HKjYp72RUXbLbJ5KwqKMtZx1Ku43K1nf46VUUKdz
2tZs+/qVE9TxntzhTxor6Zon6T1EBiA9wAZKBIj3XQq5JPcbakqCW2C9Hbp8zeGR
dHWHbVZgEdPK7oMlROKZBB7f09+7kR+Igf0lxDj8reyqA6xf0lEY3ADlIyxyllcR
KZ52LDZA5ZfGn4vDchrjNmL3zUwTD36P8/s8sO86bBR6HqaQd33nLfJ8pWeQBlCA
aLVlfdkFUQM3FZSrAd4V9y5wIAIuq0TCEO8rGMER34Q8SmdEpeEprKgbRSP+Ypul
klNp8VJOIZe4yzQdzcG9jGD40lkjbzgzPSioA1KrHRo8LOTY6htvDCCvqNmgkBvl
H9W1nLm63ojZ9cEb54/N+dV0MiwdjU/K4WdD+30yXuufNSTbPp1KFbijA6FWwMf2
5sZm5219Uv9q+iglm5Fn8OI22LhP0RyfZYhxcFyJARcfBNaJc7P2lLQ+btd5JALb
4tiineuyNLKAKS942h8ggoavrXhIpEtoEXXRIzSXxA4UA6lRChZJAqRVkIuzM/a6
uoSMYXmsqXblJMsW00go21N26wGkQszuNgYHve6S+F+ZHrfl4GixspGhFkjaSXcf
hUb2Wx4Ycr5IChRTYOVjw3eOdlDb0hFPMxuTbhW6/acKjgxr/Am56cAT+CAEIByq
iV1sZyOSIdBVntRTttctpCjSjMOUWCKdOOUU/LKxIED5AvHVrC5Ya7MD4wHpfweL
Ee/enPHxvcymS7GduMpP+hfy1VK7XEw13aOmuG5A+MLh/bG1dp+BFmOBPz4eekpQ
rGle63zQymw7y0s9GGv+QD1GAXHlwNmFVIMacVZ2Kt9DKFMA7GKLATcrPvMbieJ3
xVn2MljPeymbpsga0yKsJ26YAgY4vsBkS24DARzsuS7OGlrZW7Dew00i7HEEEuXE
/qcOi4Mzj/NMsUKITYgqfL8PasRwoQen644GSPMRO2lELBfYMwaYKubqVGE9UoUI
j8rMCcXz82dE/nwy2FRiKuomc2c/8WknW15jfbTIvUOyo+C/ccj3GnTFHRgryFkJ
jCliQUIeeMsuABHujSIh0IMaq276/IOcpO65XQ+WXztL/t/1xmtF1CZmo4DiaGCA
f/59SXt5jaZ8GTF+Pzhk54PK2JLV/rL01dtQb0NDdsbID4OuX9XU27oPR8icPLUp
mMrar8knxL8FBeF6q16k40Qtc2yHysqy9arOIIHBtlCWIO+gs/RAinHMzc335oJU
Mx5wOLa0aVxRNMFkofw1er7vZw8N+krq0wNqNDMQjNrTK+I9oBiLgUe5jLdq8orQ
/H+GT3wU+8z3OWoAr3hPAHbrj9hwIY1UfwGeM+zk765j3d3Xvs/xmSi4PLORElid
noAne3HIaK5p0x4HESYRojJ5UNwTijR75H/Uw1ctOYymItbiimhPGXXJcfvJ9KE/
AbO7EPXgTbTyZvGKdSg2FUIuHgDgdmbiQk6gfY2NLBW2oi1ZVGz0BnrEChVkQdY+
1lQCFj7D7CchADCbFEGzL3yqOSU02ek7Y9RwB5cGoUKupl+8tgkANeRK4OtqJ+83
4WWMmHMA3F0F5ir3bgjEyiSAEj/bOkZe37Bk3Pim+UBOZHFmtOs6If27jOxjB68P
5DMw3AAMQ/W5FNulKgx94MN3NZ5bZXkzaaefD8VfwdHtLghj7ypBmHITkOFLjOab
Jc0yV6sRMlpxeSLM9dxTsvpS74XpZA3vhAkW5tJ69XZWqgEPRScNMkMh9yqHnAMR
4tfXpDquIfxJ8eMR3B69MC4uEsWbjQN3qOYQrO7dCG6Nkbw9DDr/fx3Z4yKtCfCG
7JMPEPA/qqL7Fg8V0g6BJSOsWOsvig6E6fHtze7lnbbHfXKYtzj4Ov0k02um/uza
Fg1+Y3OWU3Kdwd+2GRk3xgAUTGuchHslPe6WEGkglhy8JJTHscHN1IuYW2Ksbdiy
HF8YP7w2aQq4F6acTgt+DwXID9Bx/FZcIYdQBmGuI/hECvlf309CxUonoPfx9K5c
sh9kiSifC3ACv4qimI+j8TMDIniRp1kwMpG6OVcVdmwcImWXSDcMJokg33Yj9SVM
XnEhjIeEFkIYUsBxBQBgojJBuiyHYw44aqDPohowlFyP+wCS37TA/b0uhyY16VQH
9RQ8mOC1bC++pPQTm5WbMV3O+R5s7G024F9gGwKMct4NnGg9lf8Z4N4AXYX7lwST
XzwWsTOXxBoBr980OSrkzjkF38xL7pex7Y+sdV4e4lZw9j2YtU9veuOgaCAgs+FL
4HhMhNah7Z4ho4sYZqNIBWejf/dXIMMg4K9YaToyDS3qu8wOVu4UNgDZ8XqVdRYR
b3+da+peKpIYaevNpLyOW22JGd28cTRK14/nJrWHbqpHuq7YZTayslRmbe3UiRbs
N3j0+By30x9C0My3/Ri1820PgxP8zPY8oiZdubslbZv7/dHEDh9wsiinahrTdb+t
1Uh2C09edBSvKsCtrLcET8lOZtL4k4ma4VdAVK15sLzEbaWQ9/XtuB2VhmkO9TFl
AylIvsYXHHA/z0fHb5xzkVdZZ9DIS045KRnw5ZfjkNmMDvOZeD/TUh1brFTWLgCI
Ap5OZWmEb8MJLETKucUF+SxeD+DjLSpjE0qUNz2AjkiQuz98OLNonEZqavW1mtUU
GqE5dlUYQgb621F36M+QereTStoyfsanGRKfszpK0RMJMomFWly8Z14ASdsX6CGi
VhkDxh+RnCobioGLFsXvHYZzNRDTS+cb2zxhgnIpEkoLAj2WUhBmn3FUaVdWdz6H
CD+u/nnMckN+RrTrXfK5nNecHfakT081A8xdtRx5T4nivRwT8bYsHlQUe/eNz+Oh
ezkM874WgIylzJtLlt5vgDfPc+gU4o8IU0gAXyaCgkStBjS2wBpxV6C3LY1qSF10
9yhw6CbHCQU1GTJAEZmWw12fDS2ST9gFp7bzaPI2FMpYI7NHGOOuBbe4wkgu2Psu
ga/U9tBQSi46Bs+qz9atbYJvEubkf/RX1TVpmNOzkbwInwszlSx3Plx5S6SKozxf
HH+UC1VFY3RBQN4b8QaG28IqaFsnlv95Tj4h+e8BDM8JhZo1AD+hrwIU4BzFFm7R
hwfwvXRzjs7mHRinm8oqcERmz7OUkLMVOzEEeYHFMNo0TvZb/V6J3Fz+acQ5N3hy
Rx8i+Id1FHibmTtVKRnR4JCJiFsF54+wTt1KnkaIQ9uCn8vvBqfbZMzy+WbSMs2j
2aGtxPUfUQtrK+7VPf22aQdf0ati07zVkmaLolL/dx0Gx5AeJT6znnYe98vLJrFx
9rAEmOPhAsT/4nxahq5XfzWHAU9SLaAVii4a77LUcfH30ylatXixILy9+1oLasSs
HPeahFKeGmJDkzrgGkLjrR2c0HpPUFFe5T8+jEbXcKXLuuoK3vDR9eIVT9tQLHLV
91vDBQYTx+PBoMPLV5WsRZdosqTavk9PC8GEH/R4GCBx++1ljFGU398tCo8BiqGK
52RofXP60r5rtdKf12dKO3PENYkArBN9CzgTIvNBPzj2fiEdGhPwaa0oVwzZ/pzi
Th4/sztuu0RDjUeVB6DlFS3s1IylokLqg6YIlLMYonoBHKugyICy6bat0IOb6Kvj
nXOy+qrGao9iQQUIcG6/vp06I2e3vmE3RwgKKTtoFiwNOVGB6i2YUsMZQ0frS53g
SdbZrJAY2tUC3ba34A3DinlKSWbY1CW83OySAXjbPU/oR0+YFPDMA82DHiaZAs6c
EzrxQ5mA1sSAsBizXxTaIEQP3ummwD2pbxRDlkI0lj9jE71Hsci6MEBf8eVfL0kg
S/O+Yp8hBeLxS+f2VImQ0GnbjcR2ijhxKaXf5ka+z4dkfsBZ5Y81AYHuvgNrz3DR
IAPAeJs5tgeooldi2Pt2xOQLi1xijS4Rs30voZ0Lc5uTl/pbqDndLHNGikVu85Z4
gbQEdmSD+HuyDa24BhuoYVIcNOL7VtMY4E9aIes+k1aFgnYwSKedT8wfBkqaFBwx
tv93YmKWV/PcKRPVE59p2z1av6pn8qeZyF+48t9MuUyAqpjaKTvmT4tT1SWqcR9F
xcjcICLbsm92yzfwfby9IU9urt+aft5JBANw1q4re/NlGIWnTy0HfLO1l/33RR1s
E/7Q9tR0Oe+o/9ku38svUcZ8ebL8iz2ySgnm/zq0aS+hrhGMCiENwlqIYK/nyFv2
7E6Lu8yfkfh03X2NmVxrOnQHkZeh3pw7Us/DETx0TCUGhnbxbgEFnqUXbg0x/asV
bS97UHFLe24O+sl4L1/rZaxhQWSai6f4WhPhHs7LXLsZ+ot0ijk1OsQfhBuPFswk
d2mhUXBb997mwA4tLkcf97L8VR7uor8c/pWCkSf5Z6cy7aFM6vwtsmYJvGwioeaE
206HjqArjsFQI73HGKr8azbQlZAJErbwb2xL7VLgPDpGQPS4YSVQ4Vsja42iaq35
4LbIGTAcYHGxWdMDVXYh0UBEOA3RtFwNwbTBAkzZB71QGAehzcIiunDYatU1ufSW
IaSTkXcL8EUhg4Pe08ZFaDHnSzq1HJSbovg/AN4cq9TiWVD80YHOzjY5KfiNn3aS
3PtVkKQy8PsxxEpbMjcBTuB3B8xHMOE1YRuKVEdsCRBqd+vHouKlQNN9IQ7nt0bV
Co3fZSWuVzavHk5uTcSBNno6itThbEzwPbpKzaUH92Hu52dZrDzRFES1/Aj/ih0U
tYLGfdtje3fmFtspLouesVSZc2/ovXeJob26A6ey0ZY96kQZKGGt/V1jyabiqpGm
gwll4GLo7LVNmr7E7e2oM4h7d2dvW0rTWR1F7KDQvTZcNcpqr3InHr7UjNsGrDYl
q/cjhBsD02SVfCQRgNkY08A4Od/BM4W1/4Gj2aqW91gZENOo0JHpYImjPcZ1qHbS
hkTGJ6+ll9oN2RUEjem8l8Yx3Xz94YBTu6g+9HwFXmM+DoJVhy+1JUr23YhTfWJi
2VRYMKleucGIVs9Jt4uXa1CFQQ9qUzwudRG41Jfi1w92aQbrI+GloG8/9fdK8aN2
eG5sRiULSlsitoHR4XwHSsh63+zQakAk+GqhPI3pOZRqLT2jNkhSnI31kLsMhiOJ
K9328E6m8Lb4DIOEVLPxkcMHVCaCq2u88t8gFv/NgCDW8+DVWkjRMh/8hXxaUr9W
u01euaZI3UEUvaNJIrBs+WxJOKdh3MTWiDszCn1rsDpgs65Pzb2ALlE+c/gEzDNa
vJ60/6JT7n7f53kcYo8ZToz/FGBp1VF40XuwqyPv+Dt9jhL9S3UFDinAUaoPUXjy
rJ1FBMBlDsEgHcuXW1M0aRW5cmonrNZUhKzholZ65kVzQfFZLJkrtVlphcaNB5CY
hYKHl3vUUZi8M6SzCWHZAqpt4mCjy8Q7oInPuA6Q6uDg4m7pzL6hXVhxJVgY8Oan
yb8EBRvzTxXPCULk2TiRlyH49AxX4DD8gT8WJpVbNL9LE53LopcAo7+KlDcv1dEK
wTI6UMjTtWIlc1SMy84kol98uz7tUx2oxnr98cJw4MM7Kf4AibiuoU0ZwYEaknBY
cWlGwta6zj4A/Z0DkLVv+2qjW0ntF1zJDXz0yBi/tjCE0E4uoGoWetPVSIL+WyB8
isCJDHgejW2xE4CBefwU450fqtCdZ3nknf2vwvNmvwHSzuXtcVeQJXuKj2EyL+9g
yACoE64r73i8pRJ3gHdSC96AQL7s+2y64dXKyeiG1l6G3uAeLrdCUjkWjTsUggfB
dLWsn1x0gd609IUB/w651ZqPAwKf/21s84jxDQKEkC5lXo6GYQuzmVDSeYNGuAKd
Txyw5BjgmkF4ndJlnEzAanpEi9BnClKl5WVqRu6ecl+Yz6r3n5ApEqq1fJNC8Iwi
urVoqNFZVSuqPF7pligDkJ/1cV6EtDkUNo1yqCgKic1RaopII3+t2IK5DPxI4Etv
Ec6XhLmrkUeA0OGgIuJL8niKtQnxvGJzyHc+9IUkDGIBtFgTyww2xutQVUpY1hDy
EIiOOtCFODRXHYcXvQLrmdJKGQZ4ECOdvwSz8hbgW2WgnkIz0vGvwwq8uEsm26bc
6frIVzYbXOKwLt4Ru4lvEJbJOxmwB4XmR8X5XVFxFhXOIV7ZtG/4oj6cMDrwrkQu
+lTU/jBAG0Dw3hLw4S0AzMa3dRpeHByaqMKbPBpUqTqxG5h0+aaCyUgX1R4t/yAD
HBfO6d0waBGeiNeVqXlwQRTlIZ3hDy7OSMUxQ71V3SEsVlT3dhloOGDo1RZuNvT6
SecT8sOQzWhQbB8LZ3DN4E5sP1y4X+E5LhT+WkKnFocA4VZLCvZHAkd0jjlKlb/W
NI1QB2hpU8hRhjXZ4rXoeTgCP9G8WI3+xnAaxVJ7Gz8wfjCak6OaAWlnR6QfwhX+
72fJPlx0JK42t0oDcTgO50u2/52qR+arvpoWo/5vvqdH7chHXTyKk2sIohk26RMb
xsi/vCH1MOVYY5jvt1rarC3pRLVgwatLNlY9+qYbgkSPVYaHes/j7Z6Qmr1xIkH0
RgVh2va+njywANFba10xnj1w7bG1fA9e6nGwfLUH9ETXrnfJZm788IyeNYhzMCip
wQYNfVO4t0YVWyxy8Nn4LB5XQx8ffy6NwEA0X7C5MUQI815N3XVjZ3Lebo9MdGMg
Huh85GmvkT+33SJ47767qUbzERUtylp6M9XaD+xMrPl07fu+FQQK3aamAAD4AkI7
nCqCt5eLvs8SqkmuY+TE2XjvPK+8v82pGr5oVDJhGNESCb/DZYOJFFF/eF/a2Q9G
0+9LT9ujxJDw79qrtvvQn/HU8ueq5IOzxc2fL1pGD7gVs1jQWUoEzaE7wiu9ST7c
S6oj2U/+/U/EkK88Liqa1qpGCeNN/3jMEwMa+7eNg1YK8P4D/I33NF7VaxjH3Liy
xXGpmhVEiOITt8YKeHxnjmIxa6wDaq7iNQrJB1BGAARnBcmIzfJob7PiC8UYmhGB
KQ4Jr7vsyHKElgtAXsll5VLT8194MJ+/wCxHaC7vy1Z1P8IKgEsIHF5VZfSkj7vj
Ovyglj0XncDoQ9eKG3faiwjJ6eDrJ1T9XvtGNDE7ehvdgpTnJ5KDrf/Eunady+qe
zWrDMJbPYQ7LCyEFNT7kMhcemNMyfw1tbTlWKzTRtFSpHmpESRBx9zYNjoww74e3
6SeLMmOigct6NnZ7+ELqEZptgqUb8e569WcHiWJ+WWVzIEI9yJJ88f52hYSHr4vh
S+WUkWgC2qEvRkXrS5H1TtUKpB60/09WSblR/5Z8m5nOQWIEgzsq2or3INCCkXB0
VfZGbjL5A1VLB/7NMILH9xkws1dLU9Nn8SvBnOsUHYtrQO5dvzdcqVfo9D2db/nY
fW8LfKaw8w/kZIk/wRzfEWd4KCJlxZP/L+dbW2xJu8mFajCpws91Y1jbJPAt9g2f
q/EiIdJTkBlwp7ft1rO7aVFHBSwwDmT09tDJXHcCXAwFiy0Xm8g+Z99Hvk+19MLX
bHQ6V/W3kk2CNCUCh1yLDKJ/0uOSDqy3UvNBaBuu2xEtAD1WREX+rNNk3/3hA7G/
2WGXJQPYipBIyn71OQckK3ouP0c4nTZTuQBSOoZepv0NndUCJnQrFUYQxSDgN1lK
ro4zlQT1+xxp5wG8+xXeIqV/NlbgYH+T0FD94gx1NH5fP1p+B/O7k72V6eIN7KZu
eLLzp93RYUIiLk9YbAf5DGgv/Vx+pPTW+jzVYpcftIYYqDHcEEPKWcF/YMa6Pqfr
ecBSHZzmkp9GVZ3eW45mNTVYobKrixD9ZK5931HqxfHJcU9x4gRWaH/Z0+aTtvjT
NfsLdHf66bzxe2bbOkRPlMUoQEVaJcJXzlOxYUFfOwweCt2n2SPY42VIpKXgtntJ
/+DE0xnj0ftjQBQDUK7Bd5BZuqLTTIto7/UeNG6tCqNyPxGAGj+cvgHVQWmZcQMn
UiOSM8p6SxGNVBixVAGuf6Q7u5VhJiC3L4qPFhphz//5EfwoVJ2IaZhkNHAEe6ZA
uaZCDQeXCrP5tim5qqkyZS05dwEkOMcE2xjNZvPAoJa/eBWPf4hPoPPHZqr6TDnO
bPuiK8KvvY0xkoaQ/p7JK8/evRD6MJsGVccz1kGsMGgeGWthFMDXZWQeMoOdVw5T
YbgFiUOnopCXwLV/lMUFFpZIHqcPwZuGZUPSeH1n7yLw5rvRnrrNPyUvyM3XEpWQ
QlPownXjXq4gWMzVvOV0+I7hSZ6gNyDXw733ckM10jnHUTvChsbONiZOX+rNpQIO
84pyQI5lGp6pUQNBUEcBFo+WO5qm7ud2nu+5AHxSMc6y5jWrdf7QJFIw6gnHtWhx
ksIyuqLS/j1Fth9zZMyKpQTrgft32Q9coXrzahPkvCXfUQvV12qX73JVZr7kyb3y
MhknGuPu7Z9UYqL3naxoY+fGe03032zxpa8NlFQs1+A6TYb4yBOCJ7hkz2aC0Iz5
0xBnkHwdiKqjbpMDlzpXjY0B0Sjp0D28XIMnzJYwPuA7hmx3QowK0Naf9pdR4ru1
9TI1cB4yvn/KYJk3xnBUiBhJzltYPMYo2NHxHRGO4hJkm+Z5DdI7l2F5oxS9Ehgp
aMsWT/IlDde9+HRvnOW5OsH61CnMJJJTyfhgCtTrZB9Z0sd4NjzGLcRBFK/IvPpn
P/CW5elZXeLQy2pghDba9xy1kFmR+jhEVJ5/o7+S0S3LbTf3HIGW0dBq2OTr/uaw
+z2UMyUlm1a2f5IN5Rl90h/roVQobibi5AYC5AF+Ecbqs1jYBdv8vMWdzINC2CFu
avNbNxmK25vLgSYPNq0LPkUK+WWSKb3aqoFMzj6XJl2VTFWuOrLyRUbpJ17cRw2M
AfYVm0yX4NT0YwKdQ5gnL4rb+YHN2O3AYy5SfhZgiTlxXa+pyWtJwuCcvD7aZhY6
rNTZ/g1oB3osHNit/I47mZ9GaKL8edGhuISYYEp3MtDLIAYe85KoMP41JCP0K8a3
eztjEhUH1nHn6vJUpw0voWnVS2DVabDxRqQpNXsmEQfhBNHoB5iVJr6QgECdtx5D
Jk0jH1BNjyIwr6vE9htZ53Hff8+uM8jVtXCmdX7jaAhTv1ZWV9lXMIraMwa0ECXC
PYx7yrvsUrCt1tJasFFDI069UjuqrJxg3/lU5fn/gfjRxutBrXZyrKL9ahwBy43Q
Xmo66S139FK5nYEb6j5JeMuX0upP6IG5EoaAiJJGXanntuIDb8IGQtgJosfN4/h2
vcRjrMtX8J6guzH7amTIhcXsxfSZMm/UZI3sQSkgx8qDd/oHIvKEz+4mx3h6Nh0Z
yjmTp0mgpVYdtm1QzVQ3uMw6QN0AAEGSOy+MlcGu+mGbWM/fKK/fSDRgo6ueu6a8
9xAyl1ePF/w3h8LIfeyLYYoswVXBxVqNXbWu9vzgvlvr5M4SrgW3V/wMglQjSmpj
BUjwMSxZ4EB7FyvQ/McD004aASPXjemnLJZndCthav26ja8OwG1owPA1DwGgsbi1
dygoGJHQEHNSVygOA7fdq2maYzTGdVtoClODBt1cebRp08YLnb/IQzC+eBN2TH7P
jD8DU+rY3pEEq5cj5poOTwd0rqeH8e/5z9sz1ilvaDsKZjUmUPYS/U6ZJVY75Prh
kN6PBbSUgO5O37zyRuPejI04Aa8N6vQ1t10RvYH/u2+pXLvtjrUgUKm40dN7uuZK
mXsb0eBeJZ+CkgRK7wf161ZFbQXzjw0+dfQGqMl6hsr5Wa84o5sRsvco/RDaIUCR
XKEJyeuN4+JHTM73wKzZQCO2zKHkMHeW0SSOiaV2BnNkiarrYEa8dVFXY5ltrx0s
V8K52witKnNabj+fHoDTN7+MVJYk1e2y9s1TDKlF2o1KpzEiTmGueKmhiddm+xCd
uw2wpRquXp9CjYLiQGVaq1dRN68Dt8uOCyRi4ID6HI56G6BbR3WXJb/Ka1yfCScR
KwR2uJw5K/w0xEb7ErICeVqcCf8ieRvoaEf74w8uXMBSuymeXRIIj+Fp6Trn1XW4
QPYIJhkIUwHk01//QWeMYiQ47HRr7SayHMGy60g2dsClfPBFV00wvVcBwX2ZpPwc
RE1PqQrXd4KJZtPn9PCyFlbmj+w3DMeDY5XAmoXyeKwyjBQUhR8JlEkhG54/M/C7
s+Bmgzfst+WswrQoriPVJPu2zwydDgRUJxmcAkCB+nNl/riUXHbGFwZBveLT7Gkl
d1mlxEqJgIZPXSKn0QkydBcINg2WjPrgGoOM+Ot4SC+g5SKwi9Fz82vstOeNP39l
sAYxLf6ehocCLy8HwBXkU4VHSb3xamzP6+wCHdIMRCIPo/JfFyY1EyIuCIpWR6mI
Y5yPl6BNEl2LD9hhl7pefNKr7aw24nxgCghqRZw0Otg9Rj9uqwWjCQTtriK0w9V6
RQzqBKGFl/lJhmShXaHnBSDmMX8WZK16QaH0MsMaEgNlAcitRkAM3i+HELLe5T4V
ULT8rm0dMaRzA1BymHZw8Hg3a3/J7VkhnPLUjpLelbSB8BGJeGPCXGeQEBHsCRIq
HA55A8FOAppKNDzpggQ7Vsc3LoqdZNqhZogfHCrEAz/AE15Hckj9evxKLhlY6+n/
GRXkp6i16u1Tu0s3c9tHBHeVz9fdCab2qN90SZox4llYJxwkxW5MR/4tfhKUxn+W
vkRjBLADk0w8NDfWUMZPFkFVHOMxdB/9rirQ8rCZmmXwwSzn4Nkv0/5SijB4aWlt
j/I/BqA01XZHWVtgeA/RzPXZA25lgux9l58OIB9Bmuv0Sh+2pPqQuOCJe7RgSfAC
TUABBDY1q0YUn82SBzprhMKPfoZSNmyaOxVAv+dRtyWjH5HTU+aeIgPIf7i3D8/k
v/fVmRhUI7BJEsH92TLEH6nAicAVcJGqRD3u5JrF+b6B2ocm5tTvKCYTpubTnJTl
TtQxEFoGOdbJ00sD3bCCUQGJ2hN3l0mBqWQKFdxRP+HcYjeDQ51JWO1LjrDeW8BL
GMnsITVmy4axqYzZjJBEMBjyw/NDyYCIgiqW6CrEqrT0PaG9ucsYcbJAFhX6g1tm
nnJ9KEjMjqVrl8pphXdduhbOYL76gYfUBqst5Vx3vuEsZpi2nRRss98XAFja13nN
0SgBD7kGd8khg7hVf/Q151voXS5iWPDI/cdJkjDkH04yHdcsEOhHFRS9HFYEWNjX
JbBVBuvUCiRvYRJ2S1SxD21F2DjjM3K+M7W6nKLv8kgkoHWWTSRU0sXA6HadEoBl
FCncdgoyrAVzmveRNZIl9XmIl/ci/+jZ5U4S0rq1ylfFO2gj0Mk7iYAnw8WxZl6x
Q/dwCjvdCAjMJkdvHewV9J23EgLIIO3b8O+HZdYBQ1H4MvwjN0lmf+EpzKN5qH1q
BoFqjew4j7aH8oR6A+nocBeLtrOibVD5XpKwf1/VQSQWu6FejBYT1gwAgOEYpTJO
LOkb1TVnZhmllIGhpROzf+CvgyushsevIYqpGTN4XQfg0DACEjQvhPvPhXWYRyke
OOOWvD2gasW5yJuLrkdkFNF3KsU0rQEGcdOJHf/8VKAWVd9mtipdrDDUhuWV7TPx
AFBodjIHqqVK5/X4J9PG5oBv+Tns6u30UdiH339kelh4U/EMGw/GKOGSMSreE/li
voOdEd7TSZlTgFaY3kvnTE+D3QPejjrKIw4AKZ0TmjdPMFAT27akF9HVYn+o/GqY
z/RHHgNXyffy6C1szr1kH8yd9b/lsq2+QB/Bdmwtl1B/QQVSE6cG3nkEJMJOse+T
dn7LW28fMKuTOh0/9UftZ+Wn8g7/8mRULgzFXAChRVAwF1eG5fUxz9MyPk2DVN15
TIfEtRZRAFRWi1EOZxGeFx+38bXA89QZxbfYc0oDQLCSyrlKL45BR16m5ZjWl8ti
1d/HyJClakfuouIJnQk725ouSG2wjLwu8TSolacjzkL57ajan7O/J0+W7DlG3sni
r14wsHFBPfLjWQn/k6Zkyo9ZcrP+gFEk14Yt0N3vWOPkB27SUh5X+/h7bQkC1wY5
J0KMiV44sRwT8031mS8Uj88hFdABfCYvaP+5cjbsS9/G/M8/KeFZskMXHADkFFfW
w9DI118nt13DSNdRP7c5Y/cnLdxcQgmvecrTHQyi0zbIJsLdowQ2s2Gt9yN0Iycm
v6C1jG9s/Maar7CMZwiSu1itmNworIAwc0RgFcN44W7yhSPFDjZ7bUp/F/YVCfmm
tYQx3bUYS/EBOgPCuwyeI5ZTIEuxbuEv7K/neBPUD0qRI3X4ONr5gulPUw1e18aI
ISbZ9WIXiH7ZcLy+QroNTaWsfbH0m7h/AjbP4wc7ym6h8ADsoOrykk3ZHKlVZAyQ
L1Npuoo5jcMYsGqgr5VfmkeIqdR9xs2t33zJ9k4wxY3u9kssMX1A37/Lhj/qu6Mf
miLXAKBcTN1nOVJqgPZR1HlnISPrmch7jz5U5jMVYw2tqm3nDcw3i8YFTXZ7Ho/C
q1ZSC/2muY5CUZUBYtQ7L2BfyvadLHbrVDXFiDeyqK2f+gQdxcrRxBcT5yqII8lw
iKXONbnT0dDD+7RAbvQWiqJukgXTlxnACGCVAVeufPffthw/PnQQ8rq1wZcmYo0I
gF6kD4MMEKP0dITXkcHB3wmi9SRGrOQfH8ZGCfCQARNsnPTa2y1fCwtBgXdMVOPD
yN7C2wWZ9d8y+zr8L7dWJevFGpvv2Dq7UZcbALHLAO5DJ2FFOV12fHp0sDkEp6Pm
nD7HCSGiciFyKVStKQrMTQFswTfyyrAMwIhjZxp2ZUJTiBVneRhZNmoOGxfjVsyY
cQco6KbrRUiFZQZIAcMG1lgd7bTx5D5LaeOrCLbgI03Ezlg1nKsC+aWTCyKFuRh3
j5P3B4AYDSxVOlhSgIgKdic4olhaa9WO9FS05/nmMq8yjyJTVkPwhv6RyPOaPNsj
UrCLzAGyJ4zmKrkCPYkl1xz4HpBslo39WF9tLuc54rxFJBHsXW/YyHoEcc/Ru5ZI
xLVLTzK40kxUDw0bxsNuwXRy/etgJeVLdlIhoRLqs/jqFqdRKQ8HiKFBc8icUbj+
6C/woRwgLEfQz8q/tB11qsrB2AWZLPQmLwc+CShoy/TUZ/DfkLOaT5i1IJpKpmQ0
4krVgF6cArmDztHr8QIhap4B6kR/qayqf4i5sAXnh6mT0MVXf3WUlTDjq4N5zrIh
kAGp1pt+9dW0yl4GYQhxfBzMndEhBLfeooEO0hzSP1WdEv5O4T8FeTtBrNuX6BP8
wWBn2CV8MQVua1JRF9TA9ns4zY4QIDX/tjzqXUjSVJE9aNYw3iIsg9/fOmYlIoyx
l3RAFXErAXLQs7BihYI1ftSxeCQg3gfAFTmEZVW6Mm1JyAGrZNiUL8r2E8ejisvq
yLzbzxzx/8SNcA8q3feg7Gztr7SupZf6EDqy4FpV97i4q682fXnMARu16JjrKJzC
fYrVYR2oWPVZmXcUW/xt+InjamJlqnvMp4pGHTwdZNYaZkr4Jt57pisXPDXESsjH
BxqWEkVsFVHAwTE5bwt2q/7/dq3YOws6omLhli6R3j5Hi4GRnY6V9YQH8uMFhpEz
eWn9UO7G9mtvpw4zL3nnDxxdz8DM6ZSMwNj5F/KIf8IXGhzWsVwYmv+o3Q539Ibr
DBtYDzlqX05DWOlH7I5wFLH7feoGzpv2y0UEbXIbtAahuOb0IEqbqHoDPRCkmDC9
LkBw7P0Sh7K/9CrQJAL5FwUbYzyfxxcV2dg+Np/ODmFnY/E9L9cOcyRAiy9xmST4
bnrgiFl4hIa/NJaxJW/Uevm/xJCDwwAY3uSUOxtoS0sgFqODVdSAwLqTaP2N0xB/
4EgUkVoOpLjXmJ11vnxWyje4T47ffuYDG9gKvh6i2I15bI8O4NDg/RaGGLviWCUu
Ma2zGK27AODJGHMbT/CzqTNohzHhWpJ192pLQfqO6ZNFRj9RJXy1sZhv009Vv2DT
sBSftDlZVAh23YSG3P3bwATJnOe+ZAzp7UybpLjwot2Bbb/y4qQeGNCFfzsg4Gas
R96Ui62XOtnrmvSJ2pDa2MpCFpVSXHd4GRhyQAH/8OiocXddPDtydaUJBcoDd2Rd
vdmcc/U+DipMhj7fBfiTjmff/yc9zCGwp3DKiz4F70CUX4RYuUTeSRfzz+qcDhTK
kDrrjd8McDcvZgPbYf87GNSIAPbDeF7DBG2M/MfrR6Lvygn9fUVp7kUFLLHoADBY
nVZDibWB7XSmSGVnYLE9mmvEQBBlWIUXjRoq/7QFrbpK1aWuWoWwZvzVKf4cK1Mu
DGv0pRFVjfql0RgIz2VLd9mpS3OKD8vJhYOn/b2kiHcXcsQmR4ZeX8+/blSpO1wU
sbY81Taaq3o88VA2KcLOvhiLedYzH6DdoQSTVsuLGtDfZfovfh3eVpi4fUw/kVVv
AbnqXKoODbmKHj/qIk0KMsAqldqE4YBqvBv0oVFLC+/+Qztdf+prJRCHGm1drGsm
6rrA5Fgoz0iTFTAX96HRde4A8V0a2M0we3QRWFjdOHAk04znAgSZTz3Y/F1sBZvC
MihiR7poo4Ksx1HLQR/sljD6HXnR7ubtpzcG+d56onKTyrYHFfPUsLJG2jpULB7V
bhHG5ogFJ9zdS1/Z4r8wrE6uW4f/nFirX2kACj1AJJNL+Ot6cFv6kCbB4lTmPSL1
1AdVhGBwnK224oFtnFqrSju2Rz/wAuMI5xyAWDj4vwgeOeHmuZVr3WJt6sOLEk46
LPFZVdSmHQHTz/3FZ97+sAmmze41+OKoSfgyfnyEoQ4SbLTIqrMKd/utLPmClsPa
TxaiLwppxqZRJt/+v3jO7ebj0iMV2Md7hUQRCs7JKqiq2hQ+5Z3x6oT7UbaP/s3k
iDC3wFICJZBl3C22KNTv4d325d0yDNFdbOBcDnvoU+Sioev84zmQ7kJYUWeVr3Zo
NbnYAPGbNl42xun0H0TXcjXJfEwQL2VxTiCJmu3G7JXjeph1bY+WGVYMGXOu4Nk+
DSQkYZTLAapUDpvF7gIMTu3U4rWhFY+NkcIPLc66QDkK8NLdX1Xt9f+Lfh9YWFfB
kyuGxjckhfFUKA0/jKAu0luLrqkpxIw7qEuN+eSaRekogfoG4PY/iuM4ipQvhHx3
iR1308F++/LL/Qgk7ectA9ipMgCg2lqcqAGlIcaCP16kqciEvsd8JWnuijy+omkF
9ZiJ8TGrnfbgSo6NupmpIdaM7nCk8Qk8P+SIdAYJ3mBPOd0SLYwN+FX1K3qqtAW/
eMNONEo82OTOo3yiuoxNMP4g+YuAoD84dwfcUC2A9NgRoT1LdpxrWyTrO7OGtzn0
m6ar1DofTUuBsqQAaCKFhdHuQoS8Ay5oYm6nCa31FjAPEWBlC7yumFDPcNAopU2/
lBVmnhZVg2Qdh+AGuMTktW4iP4UhS3EteJnsTCMtCN+aBgidx5x7ygrrEi7F3f/P
vRtcEIY5xHt4xvHIJHsMPlQe2KnCNjHoo7Ti8cfwqEfthDvAWs9BIlYYbXbOuhkO
Qx23WvmwrUqy09csY5xAn9gwmWzO1ZfbKRV06QsXFUNWIzhxF9hEp0gllg+FCyyd
FgJidlDELsU5OL9IG54LFNfzIE0OTOW1pYMBz+T5CVsrNMAovhIryuZGr3M/ngKI
Uh3hE+49xE8d6BTZM0Q/Hk+g5JlACNi93Aifb6DjULdD4r/2SOCb3wyqxtsMFgYD
ZspUvKuc3JxIH/icy3pjMRvPPSJWxZvUfgOh5OSDN4Tbw2KM3zh0cHbUc7MEmYjT
ZgHNKCRlWohxsC3kR6sHv3nNgFz5FKZfbOBoy1mIpfTZ2HBMZq2fj5uet4fm1lB9
SXJb3lZym1NPyDgIjnPGDiWynab4f4D+1yDioFgPcoz6amFvEiiwRj+7MoOmr0lK
hemxZGHhwrCUw+XHcDcFPjXEk93NeGiEobO+VVX75oxYzEXdCV+Elfm9k0fEC1lw
J50d3Hp9Vjoc1j/4nnAkf1gPNvX4jEiL3FyaU4KUaiQ+diqLF6RSEgzMkDjMy86O
LXlx+od6UiCla/4o3dUTFGbtQtHpSSMwC0PO61JpwFqwsMtlblMFe4+1kyTp+ni4
it3XsTl8/4zsMA9JzytqGPWryIaMEQBkDzMVpKHfCsh5MRobg1WS1ihxjmP+vXIM
k9bBN0V6MYFHSvQulfLHAhlmmwVPseg595dWB63f5TB6ZZz+TJSzO5mo3gF6/s49
8Zvz2ALjKD7LwD+hIXd40oY7sXxr09sbCsdgrFY4WrBGu6I6Tn6s1oItzaIuEypc
6obOwxVbc8Rbfuv9qnMzCfgjkP5gCZ5lSQRMgw0WnSWKeI15lcsK2P+AvJwr44Hv
aGANKuxDTetcRhsfZnVq0Aatm6IxdfTxmKwajr0wcPSENWUgx0oxsbyuaV2JbvAE
7E0aUy7CfEppmVMlAaMMpbgYhHWPoHPVB9JJb5G/KdbOd2lPtt44tI/UaQIEIFu3
udCjPMSs/KUwF8DWECrMpQggKi5DUiirmwR0kZV4EV5IUrmaSO3MlDPzpwKf/MW5
h2dWdo0NYsagc9BhQnWw8yp2WuAG9Xs1bVs4AK3YOa2ATz7JvV6OQHSa1CtsGOCz
FpoACcXBwlBTCxiOr3zwjaR+AA8kwPn8o0i7MwpZWPASfebIXSxaMgdjMkuRhF4w
iu2R4tmloFUktnDDCgwvESZ8DVVfo+R4pEqpLMYwXo631VeI0SkBGL6f4Z9CzUWd
HwWQMOT4dN/qscXblQJkhqn/JF4SI+FqjJ5l2Qa4N47kzZhfYh0jIkXty5EqK7Oj
AylrlmpgZYtM6eNsk6j41kVOnWPkzYmemJvHLgQKpPE38syG+ddv7Rkz0t6qjpA8
/1ao4liJrCBXkBwJro0ilyH1UT4CNyfqGXdUnAmHd/xE6Y7JYpmYA8FA3s7Ks0Dq
P3FxCMV8q3E4GRa/p+vffgCnrRzhmhozyrMY4xwL/aabmc2G4Pb1tjsjXxV5+RjF
ajcLcv3hOzT2Dqlmawo+lnfCvG6qva1VgLa8nvgA48Po1PqF/aBodD5HIC3j99YU
0+UhSO3YyFElCW4H4tumsvmt6TRFrKgL64e7BUYC4/JQwu6nivoogS5zxr8zStCn
esywnpY+v5sVKOJEh9iw4hK/ExRpx2JacD2WhK0iM+qhxncD08kjyzJr6F992P3h
YPiEo02v07vdE73v3atL8+893nmH68SpS6gnsGz998b9AQnkpGf78JjsSTSXAIcl
pS3FTc1YpGEmI+hEmRNeweToyjdchJLxzMPbYfPhuoQHvKD1fLAvb8Hg9rdy3ibO
xCIV4kZLgmkEmqt8ihVJ/PRf3h0LEVGygbI+jV4CtindeXa2NEANMroDfXR9Sk2/
EtORE1DPNW6WBPugM+UlFW1eRhGvZSg9O+cPKUUb2oU7o1nwgeSdJCPg+KNXGwWc
x7yb66JYZKn1EqMKyuvpbomNyBJ/CVgHBB2bZSdKIQEnxipIT+0D+qDohaNN29za
SdGur8NsxxpANv+gctk1KVyhLskmVMJiEQcL8f6F0cODyfor6S5BR8+ceUWpQl46
pgpA3tAOT7rYEPnc6dUI0sVHmGhxArZbFX0zVkWdeodkcn9St/Q+k5VaxBHNcz+9
tr08vT01Bxfug5ORLvPxJEgBJMyDKKLK950QlJQj4uv7Ycu9dNlRbQbMBzaUpuWh
9OlmGGWIDeIOM2kUb2C9OjlQkeJEki46GQp1aoZkrFGYjhVs4Dkt1O42RRTc6JN/
9rjah4E1N/IoVw/ONVvAb6u7Am6EQo7GGYAOZ8sKmhvP7Bp8rhEamE7JO+mRC/e6
yEPc6NT+pPof/s8tDNcGHmb1N6SxSuqkS0j9K4xI9sM4sd8JK3BGhY2pIOs+WdTk
/5lUucDobSOqgYpRwRKhyuELfZHgOJkjsoJqLx0HZmihTgINYsN18RnXSW47rYsT
mFRIe4Ugs4+IKPxkdO9LQ8HeyY4UnqEEWBc53zlCEegorDAllEtNhYV2Ad3spCDL
qZigR5KHVg6ikIkLiciswpzuPgSzFrlXlacGqHeh8AAMtDeDyVRcbbIgQvp6+nXU
lSI7wqjDq/e52TCPhH2znBpCXu+PnkwJTqHAdQtKDzihhSQJfyy0wHEdslnVCLdL
D6+OI9OUwASHZY4un0JBnV3qoQ7VXtTi/fu/Zs8YRw4AqDHzJwepwb9Iu8KEWZxk
CnZa3HUY0z/nO5wIcPXBtfWsClyeVwPbnf9fEGzyjHaeBRQcN6OuUI5aPWHnmQwI
utGjQ6qk688HmyK6MeEQLeMWJnS0OXvHAp4BdvV6Y4PnjGkIE4J6M9Uvzq0+O25W
9LQXOLmmZoEtiIwO3VC9/keVx9u1tZ7txDbTmSQwe4ESAm5OIm1Oqg9wC5JPnkh7
sKxUbNa4PGNmupdp6d2VgDJbZIG2urb3RpzpKJrlD8IKa4BQexDIYU1WglX4NM5B
BlHU9hAHl9w9UFZts/b7bUYhfRlt3kbABzl07caTEaMU+YkBUCGr/hcK8KMjQ6gx
LB8B/Q3ih2GqCk1AxGchkmIhf8XgOYaCXAWXZxo7u2iFdfYMhxlN3PP1LBx7uthU
dIUHZqSxBFzgDt2a/EOE5RtYdclvvZLmG5Ce+odXL4iFZtgZxZ55zYl36hNmh2UU
EoYIBuv5Qi10noueLm8608L7+pTVB5HnnF80yZGc1vN4jGJtm+t2FPth1W7i48LA
zpSfQsvhP6KFeEKwc0IdP+MXHGcnNWmeD56wsLTBXZQBh9tdvzlzDzcYHipZwrRU
xGilTnQ8tqsJR42FnbW+vEMXO04xkLkl/xcgUfgwXNrNEwLjvLXB3nL8Yt+2kAza
5MsjqCCJNzGZwd5MbCr+b0RfndVymtb4EHjyybZkNx9+lJgQ1dxjp8DDglKsva6v
YTdwDHYR/bcSBUeKNDh2ULrm+tXHHGVqUNKlNgviIJwa8hd/+euYq6MmeJTZD06F
bvMRtjjSCVh7Q5c/hWXIDn2zNRhFvavE0jXy2Z+RFDOo+CasF7HP2hIStoyhFiql
7zX+VJGh+MFpOnS2rZDhN/sNbB83QWEDHOefjR+K7MkQ9OzzZWVgO7s86ahrnDVW
SAc+mNTSbFUOWohGq9CzUfnVOtl0b/2bdEy+uxJVqhFtdhbgK/ytmI8C/Nrb/54w
PeJNfSN/jH0MMLE3Zui+lEeQaweNOPqxWSTLIhWKNE+ZGFy4dsi8+qRM3bhraUd1
9iA4716dcwhTPBXKqC6Bh/mFz0fsLcrOdsv52faWvnWfqfCW+WFE4yV9DMiatnvv
QcuTxycdGzw+IxnBy+N937oAcioIJYpl5nfdBPPcT/+yjFaWyONQxCDch2YwUeLp
przaw0InfuEFFI16emv0lLbxowRbH+dccgLUwANd9rLcI1lgcATxJxjUahfF2WIR
ix1qKDHFKnIR5GOg88IR6e6q8qa/Qt++E1miqtfdFcrY0+QRaO7NU7NSqTDkeAd7
bXEWLYXtWttfw2mHZ6dyAasj2p2RQM8TMwjNVyqUfR6XVF/iyEvtbWDmzLM4i43P
WbIf8SQocHSzEpkPIiL6TmtRquDSoc4M8c9cK/Pksb7Z8P0dkYGJPhox1HCjkMYT
U2ueLhO++OmKGFthM8rb8Ug4DP656WbGRb7wdvm9Vo4NkxQwSCnOYUXPm0oCW8aS
t7JbfNnX7/YuD9PFWjrzNohZyH+VGy+a41rwTKV2QJccXQ5rFEESMShIaBx46KYs
ZOQjvhJ5LyGLvL9uJj5kTdJmYQhU4vkElR8xhn5e5a2/z+v6joUsGyyxrNVOGiwH
rcin1IU+20X0N96SCZpX4oCzzCGogT0I2yyTGVRpvFTzpWscWqZYvspIyuidKSNl
ZJL+LPPmnqcc+r3HpGjwM5hC/f4ewoV2Nqhlv1OFzV5aUik2YbLkQBJu9RxXWbve
qv8phjcTI9umnZni2Rd75lcuyijXpFclrfAz2oc9R3YZaeQaIHEwYBTor9BkSWvx
XGuNPdirCTS0QxTckuULO4TRe0Mj8X3G83x39b8k7UuR09tgRaaHUDOx9V5jNBaE
EhYE86NFYFPQTnvdjGt0SCNtt2KQz0iiMmayJgJQ5t1eDHARCSTxUTG4k0kK549J
AK5eamFMq9zvufAuj7Vqb1BnBnuvL3RxQ1IIYwKbzgw8gvstX/b8CujH41u2ZREq
08HY0UaBbu8K+KGU9Mg5aXXJoEsTv6T6WLgRh6LbmIKOfdws9FHzxuVKYyKowRRu
aI7rlRqCEK+n+nrUrySBun9dEo8iomFcInMuyF9akPugM84nl0M75kCf0VFiXtef
Ooo5jsEuQQUtfN22SYfK27N1S1RqJiYQLsrkaYx+jp5aCrq5uktVG8eaXCCaB5mc
qKDZwD/gCEb52i9nclUw5V9ZyTYkC2VY9qgaAgcxWp34ni19qRreomy6CMdJWLeM
S2jwYiS5GlngOFzN7UanfkR6iWWwmy3zB5/9Dd8gPIIDzuNBq4XOJyAjYv4BqA9n
4VFyOyII5b2HZ3Me3sNVA21DDhWRu5Es6KtYmU7CYwc4VjrxEqVXQ1Tk7SPChMAu
JIIh9Y9q4BCjtD1uDG23vh6k1GYKZYwbQkCgBqBqWgmnj/YL7b8kghdZtLlu3eJ6
xsWFYzAbhWaYqznCz9vT7aZH4PKp4pzwKYax8KwysNk97SSEbpS1JPyFx0Yj3Ww5
g/p/AXVihhp1B83twl6f7DQnuYg/NIvUvou2B0OfGB0M6YzvyBldKPIgcvR3o6Yg
ccP+fg3Ak0l9twWXNQGi3r66na6IpV5qLgAlU4OW4ID+HQWFiiubQ/yFitAC4ozt
oDhoOQuOW22HYchUXdcvB41e3b5wQptTM2PW/65/x2BlQ2lQu9RJ+l8J0J9kOmUP
cdVkr3LiwUmfPTC42hfuAPmSGB7kOO5GZW10kQCzeXe1eNCo1kY2FP/Qvx82xyi1
8rYUDkKI2VWIfHjTmGiPCDTJ6SJTayL0kxljuxE2VefKSXFGQddbEuZ3d7NqKJwk
0a7qAiroFsdZof443zR7TL43qIQuvAoKO31FRfBxoQwI4qv9FxPMrYSlQeVIaU6j
V1rpq6ziRW1Sb2BrYYaaAgrtpkxilto8lfzI5cYpExRCYaBqjKpS9wzP41Dfk+6c
CDtwrTVGxNzHGbvsx6k6uhy+nHwGRig6Zs2I7B/fhpjRYjCwK5vW592S+U46wBX3
Cnauyx/bXlh9o8r1/GNekthSJasZaACd1VYGSgjjMudonuroLi8M0R/ZnStg5q9q
pzk4IEUe7hzGP8F+LrOsUOrP4lZv0OfsDzKuoiBlDVyjOa4LWfJeJ7hA4s2RnMWY
onh2A1Cn7aoYvab44zi3526zVWYSb9mkLvK8leeqvKaj6onpWIE3nZct5RtZrCvK
RiuBCfM0U+Xe0/1LemLH11W2+viIWfOrCkrYhmHQxDHP6fZEfzr8A21oS/t/CjHx
heXlmYtsWlFrD3dpoKM55YvSl6fXnIZP4twOEJOeYHCNkIQy0CXgaAR7SKkaBXil
pKjp192um2WQzJ0f+noH8ciqKnv3qL+0PNOE439qaYmKrl7/tMBmoLCUOh7T9kZx
JwXa/8gpw3FBL0O6jXEhgELtYlxuHFKoQaCgMvtes1ZN+ev6Q37oKFiDRSwpzoOC
tp/OcUS5HoE+L/qrOuWJksaTbO534iNJ8rkbwha4wkqkmrf5DOmSFM6sqB8A6np2
q19jzTT7Xhc1gns+eONZ+jYqD6m9Uf6wtYsVZEwPKJmdcAHpmJxt9sY8WyVi1ivB
jY3Pm9iJEgsX90Fwdq+9LQltErAwYkDNJwUji2IrKBA8n6Y0EzWp6H1E9VbcNJ/O
i3r6E5toSn0q92j9K0bdyKyBtxn3ut9C3gKocx9itNzZ9DOEpFsnFhglVtpn+xpY
uk5pQ7rkB+feutAculJWiFVP2eyn4QthAgfSXCsywRBzFARUDBkACMj4WkQ0jvkr
KY4yI+v3ufITLtP3DbMZOLGlMrbZ1cuKyRZknGKeFIOzAw63elidlzobpS2/hFQo
nFk0owE++hYIZJOc5HIA73ylcpwVFCAqlUQmYaAS8ROHvVgyxuMPIir/AcDHXmXC
qT7h6uzbouwCJpIWS10u9sPD+/5SymycCcGD3nRo4DyE/VSBXX4fMbZxdB0sXgkW
wK48CAQ7/+KXxAHml/QtUPHYMnFGpNeXxQDCOXiCaGHPBIv/trwi/sUgVHBrM41Y
5F2dDaO05KN1uCebI9J07NUvtW3a170XBYzynjr1mWPzs0d9JHykM4nzcbutcJCu
l9eWiEGzLiat20En3Kp8is5xph8kHaZKY0A8VygBDtVUj4VTQ7RS65kgu5H06F5Q
zgy6r2zvKpPfg83LuZAa9vk/SuJi22SngojN1JW4usMmn53mc0WBPl+iyR0NV45n
g6I7KmnLg3aKVLnaHwgKq54W0yg4pz3wN/nhQKGVBaJCQ5vAiJrpnsvKmS/aHmhf
JueLiT6xTQGWb61aAx+Qz/0XDwOyPRXuv7B22UrmZ7WwbGADZ58toIxbNMs+C4kb
3kvGxVqAoEp/sfUatxf4VoQ4AfXYvFNZRz68dUCiNzRROyG66ugsAz3/kEOfAzP3
Uzvt+3pXNrou+8TKbjF0Cc+1zx1Nkrf02IsVfP796MpB+8NbdtXXRcdUs3GWlLFa
2YSZ3xO0Z3PsjEbkGAWi8IpXudq9PjGmrqlXF2mGXbnJ7kUzvmxxqvT6tFedcvfQ
CYdU0bvpGXzN4nzbWkNljyMQIZD66IPAI0QVTl48Be+bVOlH5PqlAeK888F8nUHN
YpPMqNG2UEyOqom9GUwp2qeX74woJP6B4+jIzzU9jhH3P0WCZQ3r563TutheF0Oc
MCqCqMbbzSDnLJA5AEZZ1FncD0xiVUphktTuEuBlcMYbpnl4kyBKRVJs8KrrfW3a
rMgbdUvgrvZmp3M47I7Ae1JUVE4El/lEnqc0PT6nwmRWGosMoRKpW8Jar+ojNvZi
Ww5ZI8V8x3o+93CsbbkBbbszlk3uC59U2uBVkYBGzbMr5XG6ANgv5HGDuK/NsPKk
jKFgjiNaYtHGkqvUXRyxpeO54EyOrV5+Yk3tBcCctlNbXKZVYqPmJ9+/e4R84NHm
llCaxvFf45Qy7Xmn0xsZVKjJTkkSk7kg0omC2B2/cmx95pRYCkh7S9EdvtXTQyOc
ou3cwlKXt2fxMlRW1F8dY4K77ju7bG8Pyt0rY/HfVXZK8kKS/sjYBwS7cW1LBRcm
+5uMkVXzci8B8iC3LXKsng/oMmINiEq4paU/DBGuCiZjWYEQ4GSbkbK3yGsDWf0K
n7aOiTdJ6+JCoGmDV0Vx4+/SZTTkJiNsGANioaokpOjm0pffBAtLAMIEY01RFTsc
WJrTmvALJYbr0K0ut8DUTUeSRFsrove1FPzzGu+DzM5EhDsIyuzjp5Nu6S7OE+nl
ym52UrNxiFPHs8/WkobiN46Mhw12irQGY0Tu2ZVNL4/5CWemRleMP/gIl12oIQ04
5s6V8xTJHv35D+qqKSCq1ZUCIDHyM5pOtwODgyrqdv7x+ytHd/GnY+5GZhUfQqY0
ttOldtWrqer3omQNpoDRCZtvrz+8pxVNpvt6xfN9vPCOfAZJBIy+SuG3lTirLCYA
GOMIC0uo0tthWhq4FYlDwXU6Uz4wloCo8xhDAQu1f5ekGgS2nQeQq4gTOitbChLA
OEmFPzBwaP/+UYh9zUlkL7XDaIsdIs8TxSkTCBBsVb0GmV1c8MtRzEULrfg5kARR
rVR19FujE9mu0L5dXsjSJhdAweYk6h0pFCdyqnWa1EsHXx4NYzU6c9wksZ8MPDUL
xLTNZMpREtenwDwApwLON1Jf1tjFI7izP3mm+7HOXnpIyTXB8fLzOPzBXlwRS40F
HI5GoT6N4v7IQdsDUoyozjQCyoj78arV5MNnqmu5bk8tB4RdEaTz5VpqXAqeAoxA
7W/9MaaSMdCVj+HZvRG/7PRkSQKz/XGZPULnn2KpskR+DsXBtfi3UtvVCwjyq660
mOkaOMJ86bS8ffKsSxyEBZQcoM+0IOxQKphr6hDglLvc23dV8Keo3aNFp7XQNy1G
3ZBBTC3X01tyfdD++8fbHuj+//OXyXIbIpjcrdEvDTgUR5VUx9FB25WGgFoCD7BY
kG5wcGLemFZDa+8j/AH3rohyLTwiW3jYAqqNfl8jOGMkBPiRoyU+CR3QkOjAf6pK
ntDfplZaB0Cq8Bc7r9t5Fs154vcPq3l7tnt/qrgTZcq0bA08bcM1LV2uKHQ01ioR
X3HfZcI0iGEk+l6znaO3J3O1ON60zt5TnY7+zQvrvJDkyo0Gn8yN9SG8aZtVB2im
pUY+3lh+ZLaSHVDZ4kEa8E5ktP792W5IFgdZgL8STz1dAYPNhBqj/Tu6HO9AlvKm
8VhLdrxSHytoZ842FHAZa9O3n0bmVyjIUkLTRjTBvgvcWIWEOatq1h+60AMaHM1B
w3Bmva8f8wTs05d7FbyAknYw5H0BRBES+xkIiprpet0trafIDFQucO1ELLiBzeuR
mwSPfrVUwGw7rozPFjKsGE5KHHXJ0T/DfceION+77xUXZmeRvriozIHjIHKaaa89
KVtZZIHkpef5EF5gJijzOByWq4ADxjJVLvCOTdTw5MlnL5gm2NW2yqCtw8b/vUGy
Va8Ql2mo3gltVZbyRjm8bFwZUWyGO3zZsT/5VhasfB0OdLvO31aCuLlcX6NkBSYK
8ygp9doJIX3IdDPi1Ez2tzAtTpM2N+nngvdnPv7Qk8ZknHqyL1yMDGt3LSTUp+K5
vcbFshgfB4FyPPPnAIEgV4XQYz2bWj1uwqCD7fs0wuVcMi8Xkel7RK87roTj2juM
9tQ6yMfaouWNrJOKO792CN36fuj8wY4Qqj8BGcg56hWhiBxELgQyA69CWjzkUP+d
0UGR7kWBfmES0nOAcbTPnsKhKJb6+AqbflAWEQlytM5rgzh+nEjQbqNbJELM8/+S
3jLkwOoG54hbuWBGTwSWbiln09QYKItiXOX14hW7ydQjNQZvCXTQE2jct8pQmMN5
qDaK58DLCPGAN1Dc9UrsqCNFHeX4dxq3fcxCVFdeBnYE+8xdiHtDSG5KzVvV7h+s
oJ+/Anf4EcrB+LXy/kWO3+x3p9D2TkWqiE1v91kPTAjDGFx3rXooiCgwRL/xzNs9
g9L89suE3Ar8W3Gogp7m1HmmnPI2F4PjD8ajLXd1iPOS4JpLELPcQIvYHX8Il4b0
5NDEShND1x9Poo2bxdYXAmzy1ogeZ6Bk0WnEdLjWB0Nc0kUYM6aL3StyH1bylEeW
Un0+3mki/91mVvXsEJWM8Iq0IaG5Q9eXOxZJf3OH44w+iaIzC98ZFToM+GqVZxWt
8PPEJp/nGzA7YIkMkIvKxf0wuUaO2Id/1SgWv7zZvYsDajURzri+ptpTgOsVnQ7H
vX9WAoCnUASH/+TQoRxFH8BMSoREncVTxYIqXKtafcGLssjyNj6P9t4u7hBBzeP3
nA+R3bEAl5q2QqHnKlAiHvYe0WinYDUGupio0hlzXMjFmAHYdVECNRMaIQWdRdlg
NNN5A6Svw/05mAvmrmVVN6hCPnxa0NnTXCgOWMjLWlP+cm4Mvykh6OAwscoLr/so
wNhAistj9mhfoon3XeJYsaA+yDIEsApP+93DnZ4T6/hpwv9OFLDdqOMoP0v4dAK1
L6s6d2dxEc5wXgB3l9QpU+L3YHja0U5FjeUDEeQiUX7zcmwZFI0/PaXByklQ0wkQ
Jo9s5G0Y/9LY7QjY2qrczhncoyIKuPeUBnKV4FyO4Z80CBesfy880qx+LpcLy3P8
t3nVQoPPV7OMXhoaSaWCd/Btw8g5Mt8Wqw7vu7uOszjZ9nJzFiQWOZORgJsO/UON
TbzD/HrZ5/CkSlrSe7+Cpo/khZYy1j4szF6biU7a9dCASSpsLpIBnhMnmsJbuGE4
KMIVBGHNRqZVosqPCSdUFr7TkkUZRIosRKzibnEkrhz5IZtG2YqpNdsjlle/UmWi
thBnAdch9MaIbHSIsHHUGcMq3dpzKYKdLEEVBBSwrXnUNMzXi82rc9wAOZAdohLM
tZozpm0ry1G/RbMRnGgo2Z0DMY8y5ewCMm+5J2J9kyB5+HCzHD0++0kapP8ZN86J
O7YulgegzKNgixThbsKUzPiPtO8qjdsFwJh+sE9W+9ZYTI7t7fgBGF9qzCg8pt0+
ufvwwLU1sQM/Hb6SdtMq9x10pomod6PzgWJIgyJmixahyM88q9lXIu4JmhLWB8lb
1juFPWm89p4H/b7K2Li1T9RQO/rd/z8F3etb2Qw5N/KVfA97usi2gw/o03LpszEo
/twABeQHulAPL4lWB+AedYRm/v5RodVUzLGqgDbySAfKF4IoctogR/1PbzM2hGCk
8YnHlM1ZaQBUgdFA3n2YAAzv+3zydCnAZ6SwVVdtJVVpS4fhSz3n2uYlL+ybfsLt
btGRDtM3FNC8KBwPqnUXZ4h4OZNCtODmKM2AD/eOcDSsEHaJfLPK+sqGymNiwZZ+
U05CS2FhOE4Ue2+5axq/D9UrWJOv3tK3boovlzveiNM/pUy280zDHHSVcLCESM9Z
JvJ2nbqx8pDzVs0L7Z+G0wHjB7HiDODtd9NavaGrUk9xMqZY6qK7grsk3pGYuupr
7+zd8FZSScj1Z7Y5JoAQ/TNXXKyvNl7F/WmEpEbBC0BBRfIH00L9gu82CqGBMjNd
5rL5QwzrgaiFnCH99TicSmQO8zdbxTXcM+KF7sKNRt/yz/Gd37sHO9/oHhlIjHzH
4vvx3eWF08qpCvzjTZchoFEsAd+lqZIYUQV1fkeLVQU37GU29Bri9aguPP1kq5U2
4dkTdCP2wmXfadFNTWg/+xWTCRtf3mp45WnZhqzpQFJ2T/RrlTQrixkrIEM6km+3
xoJsRzGkEMT0sTdNxfvl6F2KpRxOZwRe9fXn0ol92vi0oW8F3861NLZLUOrwZE3L
qK6tcYg9NnOJu9ZTSIvTPdnccRIHVD9qihgoYTa3JXGOomQ5PD2SN8aBZS2iJnG4
ts2pA10V9fUlzAGr2ahqXlLqHtXwA2tdrQmQkogVESuuMJ+uRGbSSmnhD8qMa2FG
wJNZ84QKU4ubp4jSSoJmtzxC2ROn+GAiovfV2Mz6/2TPb2yTLOSJvEPc7gm+UlfD
+L5MmIMcEG/6MVoH3jmGwdCESxUhon2grWoJ14Ro9x6p4qTSisbg4WTfzvzRbts9
SDmrWwOWoLdOGx6oJxCNDf1YLg1en0mYkO7K4MJoRH/4WjjpE92bl74Yp4U/N0dJ
rpjd7LaMZoBISMkIbv3U/781JrnvqVj4VhvW2tGrZgvM2LKIFRBI6Tx1f6DkAAZH
Ia+BDqeNqSIFd9AlMCCTwfGXL4Z3fQMJGhQUO+5hbHTxJC9vdI6ayDuOiK2shzGf
NmHtt81ZLeWr/eFdzlTGo6gM2Lt6oM/c5MS500mMcRcQYCOT5Pejor2ufVsiyZh6
LqtSkt9btKJJz0yZBerssYO9hsF08MeE7UjkLgKAFua+GGy+nDPbiqt5UUrMIMLU
qcbd2G4snOQGp6/J4T+z9pwLE/OXa3dGZ56jpfNwTrmx3ZI4ckPAbhHj1AMys0XA
eHzzIkaJVDb7kMeQC3WLLzKyhlfeI8fV2Qp4iuKWk939gzyLVKsBAOBvvalO+tXu
A0lvlXYkPs6UT+xNjcZ+7lZjvQbsSAM1ui7KkaRl1kFpynx81U3nQ/cRCBCp4V2Z
mlDyqcp0EbcBF0ZE5zQJkEeYtsDn821h4ADrs1e4TKNn+J/1OT8qo6bblkxHXd2p
zc0+IA/j9VUrF2PfoJK0dbEkQN/HXQsiIdHXf2E/1l7OrqVuyBNsPzjL4eAa0aQ3
aoBWIT3Q8nb0VlZXAj+J8wMzUKVGDmqiIsHcW2ex+q3mkqOqzY5yhouNEdBeClyl
n7Tmk0seiXFZbkrMjzzTVNZsG2fvkjGCHCpHTLJESM/PgtIAbnmacl2t+M3VvFEv
grW8eHIXY7zdm0Z4VFw6TkAYJV9TXFvXocbWGHoyN2nvKaHtVgBJtPTDNXikZHb3
4aldXaw8M2gRI3hqdRS+Lv2PshphtkFAz0KSu5zBjXJ8JDKRpe1yK5FWoInTjw2Y
+Pk1Bqc0IpBXBFaYUie6va+dMJgq2E2PpJMKFLAXS5QiQK6Jbl5bodgP5ZzxEdzP
FagPxXBE6FrqQuf8wn3Y8oBr+xdfakON8DGRwBg9EiNeagAWKueq8lrhA0PEilXP
QpAvumHnTGxYOOni58Ffj8PbjFKDYeSUmbvFMHsGHHx02LUQgG1E9/e74wQSYfB4
l3TZdA70A9PSzG5/6gzZjE3KiT/Nm/2DiseCtvtDVM1NlFB8MWGleM9+8dfR/B3S
79yjK0WbtRsWDcw39J/Mg/e2YLM2S4HiR/EgrEJDDdSSlcvoUnfW7nmR2mWh/V7w
K2cVMeIqCmLWlP9GfSEcu0TSpBxi5MFG0zdEDcYCsCTr2FXOK5NWnzib51nXPQTb
1ShX41qtaIXHzp4TiEw2N76lIWr7X6xrUMag/R+KJo0EJp9CUDOQ3loe759jmETd
qKnQXW2XcrZ+cWZznxNpIikohef2oDaHPdOTm9NZY7ArechwOiiVKKB5hc5isw/j
g5T9QtdRI5VISxzpNKRQ80AbjQJah/kaxmvm+bNkyDFLCVJfcZx1THCzzWRW9QZa
KjKmfP9LQvTCGwfeeonPHPQ+cyKhfJUSRDcIug5R63jqvnDC6DqrOcnyN5AopafL
ki030E11xRTnXNvY7QgzIaP0M0mMiU6Og0rKd6vWrBbma6/b/RUjbWVoeegkbmW9
wFNOZPTTb22uQU/GLpHKrL1xQz69ryNfg3NDqBtLbwhVnPdOqQrxZJmaFbAOTNL/
5qpCyqRQzAuo0TxTJ0ECW+l7CckFCc/r9fe5X5fjtwl4v1c0wfPjTncTQaill0fr
kFBS9UPK8afUW922o7DaGV8ujBCxD5STgBwvpcVjg51/3/WDdMWpWr2WvEMkHUfU
lKxhDyoUc6NML75dNF8vqSahpwC+Bm76/twXh36csbh5m3UHTJzex/fSJBQ8nfQX
c2o/SQ32JOYr7uKHMzUmo+Jx2VdM5tivL+knZnUWonBfYSYRQPARjZjt0dRIoYkS
Top6EPYgZDjStsEPhVxLi8u+5erVAofLO5BkZfBy2YaTayJfiERdray9rhOcORnD
s20+Zua8JlLOoD7I3LNZeVNvvdIU4XufRuBseYHvko4Gxhl5e+Fpe9p+MPtbK5TY
Mu/Xh4B3YDcBza6CB9JE64ZJUeZXkhf5eMhu8MFyqZCYZ2tdxV7KMn7+T1Z8Gh3o
5xgpiyhRdIG32NMU5FHITpD1oV+UmnZRCHJx6Xue7p4S/GcznUIp4mmWFEfntDOk
5qEsDdGgdX8XoNXdrDRa/XPcK5mPxm6xaB67jAOZfyYpMMQjsZWUYXX6jkZo1MVZ
86jpHmNjNnfgv33f7bmFY6DienYxcBOzEggmJfZoys2RqqiMKvfBLWCc//mXQAEW
wmbLUmreM9ujRIY2fSQFRY3+FGwMOWC99k8lFKM5IHrxwqGkhjf4bN4GsW7TZUjG
k0Suy3CFl6zuZfi5PNYXBTfSiAIHLgNRik2HDkoVg8s2glAYIFUofvwsa3QL3wSf
9ZEEkFiuZ91EbtlJZgxYOi5yHDhkMzKiUCzssuNYSSSRHuALA8mLEnS5203tJQUl
5KzvtidXXfZUL5p7nw9VJg4343IXYnhpWYp71w5pZyFd5bMKwn8jgD44DJkBfuuQ
fa4WUOKrWosEcYPJSSqjWaSWT6HdI0VyLKwZE6Rx239ybm5g34IKPMU4LT/V9Wp1
bBTJCBJyIV9NDIJ2lB0KzBZcDYTvCPmYpfj79YlIh34KvQ49Z/9+djqEQOZhuuGZ
+2XnvIjDX578YybfUjabh+31fUNxkptCjb/U9eYpR4LM0OiOOPIxbXhac/dT6oBR
rLh+8G4xlN+jeRK4muKKeRZswQdxajQNSihHWYZ0ZAnwYdfOAHvuuoair0dYtoRV
kUZTaIGh/N8xV2c3sQNEaeCt9qEVQa7BU0ZaHorp3soqfwHFjqnSRSKToi8T7APR
xODId9HZ4jdJTNIrIjipIRj7lH2czlmRT6q489TGyGVDsKM7VC5J0jGZHXhiPJ/9
x2vP67Fr/+laEbusNGBnqWCl/XQlDc50p704ubxSr26rt7Lw01XgBUz7c+W9mA9g
RFZB/pKMco9nl2jkFXa9356rkyC7juXOgLT8AqfO+66rfEDBwq+jL6P252grNFz0
a/2r9FuBvaq+pF13Z9tQ5KDtqrxTpUk34184f75D2UmEDLys6F458+sxgTs00fCr
QLpwPV5bTanGvqA2Kfw30sOVQBLESZgz/GIprBVJQS/kxz/vS9wLRt72zGIbtcZ6
1q+uMOCZRckQtyrXz431C4oPMqFYjNtdv5Wwd7pREzToUWNa5AbKIin/iRhZxbL7
jBHFZ+lO0XmLMuiZCbrJaYQy23hX9eBUMdXx0F1XYOtxuVI7sdV1BNvaOVI4RVZu
EeeIzBbQ2zJmnwWpFvIYkd87a3wtk5U5JpoFRYKCYPklz3h+43wku8xfjhmp6/EG
BcUJq7azaTRmocDB0zaJHHVVyA7bn29yvQ1ZCOkSmxMdt7lAz1ffvdoc6dmZlXUx
BAJ7sTn1E2woTx9862rY+kLzyfkd54rbpKQYV/Oy2Oeg0MNGQXkLpT6WBcHGhI/3
z/sBIflcidxPxCi2E9tm52FhJdyFPQsIIafEQIlke5FdvGiHLg+ToS4XQVtYd3MS
Sv4wLR7b8isCysHDdRNB6/Dj2o9AHZyc0At1XV3kXDDnuMY3SGtjNGeZQixXturn
RSKlv25lxXfhQktWxU26sCNlpfXHElAIPynUrKzOWj45ORy1Qxm7aoTaJjGktVK0
FYyMXDcDWNnuTNozpP6aAiaLEjHOxY7NkuIpcfAOdd2JEHbqN33qlGaEUIOq4RA0
6Z4CfWaw+eG9eLwu03kUWiCveShwr1YmtGUBATPnKuqnx95JWkCZKjXmtfH/sA2B
YPt2jptQKGoMmH+UyO7lq0rJfc4tKe9fJTAwDH7hBuBgsS/YANhb4f5UdbDU9gpE
1jLw1CTqUYLOPO+T6XAQ+OhXA3pkb/qtJKKtqe9e/wu/c7t65T09We3K3x6g2cxX
VoLZaLf8VY6VlDKSbaV45Xe9nJV9CcjKg41g/XZzpPohsK6LV0eozrjQ/hheZmb/
k3Su0ng57Uv7isWPt7JSr7B4swX0e3p65Y86xgioCoKPFDjv53cbnw6bh5IEAUMt
y0+wO2jIXGJOSTN7dzKqt1bCpNpWkj8BDDyG+F6x4sRtHkipOaV9SyzHP9vtLQxh
fTIyUYhz9LD05wEjUy+elWCw+/2SITbfkyeBU2lRc+2t0m/QsRR+MY03fyu2oi9X
jWFSHi6Ws+JUwxoDNJQnJ7RXRHrrHLxn4N2gVehJmAi3e5OPWTwj5bZ4pb58Mes7
hr2olG5mfB984dYiYR6QTovqpj748x/PeN36c/C4mmt7iDm7l5rnhAnfZqHFQqiJ
A27VqnjGcRisRZUmP7fHcpScOGQ1e4Uu5nlgPXz3Fwc0lemfJD0SazJ6BJKCta0i
Itfhu0GJRpbATeAh007DOQVKr+wtAINisL2CXGxMGGMSjE2ANjrNgAhuddzTWLUt
XJ63sBPC7vhMG14Ec546gClEmTuXs7xn2Z2Hqx4kyQIyBEV26Z9pmjGdr22So0t3
TOHgZ+BOkBqH65K9x5dTCRv3vrgot0wD+PY0ZQZFSz8Cj/5rdcenQ03JsZkoKqyF
zygVs8S5ZxCZfsYGFNcszBl0zrwLcgLqXY6HpINc4GVryt8tUSEurlTQCuDlFsTp
CyVj8DhVPyzB0o2XSoXpwByOXYDLfN29wU1MIMwWMz8gTLajDcPYLGCeMY12zC/D
V6v5ihjutJ+4qMyVYRTaVObdYy/4c2j0DrMInV/hbqBLSNzHt3pq7VU8UeW0thyW
DVdDdAwKNc6kfqJJCVSSt2m+KW2v7KPE0mPX+2jpt9xxrHcrk7F4q2vGiHnE9kaG
hHTKKgvNb7PwSqOhH8frl1s2k9qeUJlvkzeg9I7gMUJOv9bHVVLNtoFoN8VLk6aC
mbGM1ZiKJAV25hlRj0DASsyNnbkJnFAHih8vTJlUuC6YNDULWUHRozjoVGo9lK5K
8e3+EClw3oYzGoZNIAZfjT1Mez1dtkFPz5VBaYIiBSJ9x9s5tLO5hxl3dh0ZQF41
fwN5uz/whdOSw9MIUEYBHbA1ufTyfDFm6ccjKwyYJXzJxWOAqHH3m8l9ARhwC/QH
1yUQCaH9XQbCs06TZ10hc9snS5L4+DPQYamfcnesA0XGqPfufEIXEJX5HEZUVRd0
bmoGxYHSc9hUib2ehak+2133bwuCWaG9OBoB78GLSFnvYF3VuZjQl9uGbIVkDMra
A6D2vHvQlCLo1z1rhTHUrXfoukn9m4ykvQ6tsjDs2AmTRPgYb354kWadkkqZ4vRf
wfYIWIEG/+6EanxlbPK9eYuOH2VXlr5iGDHN2LfKKufP4zH+3p2u2OtR6lw9Sl7s
aeSNKQ+s+3zilu5F0MdOaLALZvNUwDC6n1czU61tTsPKs4yBGK/WirtvlGlcsEkr
GQ+i2gyiR0XpBQvLboJXL+wPL3xf28FvEiW0FaiLzPEQbWxIwnFJaSU4iRGs0AFE
ZMtbO9/Vhsmp7J6FRg33b2x402b/g6vv8PG2azl9onsmotSbbau9lhPbflJGd7ll
rihKQ67keSEOdqHPXWrJoP407wxOieFKxLgVShW6glDyuAiHFHMH8TUuy0CHMhC/
vuWQydkrh3nWaY1G4M9QTcAmUFyYp5aSefXkF4uhs+kYoFLOcuZ5Ulfpy8iQGtl2
XmXu9cpGhz1zOJP7TANZFLdgpOpcO9BricqjbyUSamSpacZBkcqiHfGfkM3mF8mE
dUjPjU+IBmsRFkJXd/io4UGaf9KjSE3/8aPPcCV5Jtede/ggJ0LsLrmZGj6K3SAI
LjUlFa1YFn196/H+yEY1gz2ds3k1NU0HsrvoArSQmiXNVlPXZwMzG2DFH8VKxGRp
dw/OEi5RNtHRCtEyqFiV5JHJil6zS43O6wAuNRhuKzAzqoKWB3IBlL2bmtVf7rRH
5EOkc2mBJ6bSKGqgp6MXJ//64qbzgpLpyg1+YnexkTzzvSwnfwW+x8AY5+B9c6VO
CnfXJrqaWqfmhcJe626SX6xdzTRU+PGpnc2uCiR+s7GhQ+p8u61QJgCd5Hzqseas
Wu3OvWf+sWaPRB2a6W5DzLiUVaggTa6/eIWdttPF9ET0JED6FbOPkr2QooSNTnsM
7PTFMx/xH8T/SuuEKjz8xNuVvgg67nE5pmTZZPKrpeECMTU+ZVsh/yro0CCd1eIg
L5kYNynYz2BK3vYPNTMROefEkwZYc1AsnDm3XZB204opL1IUOrBTOjnA5eiKlH3f
dSgpz3QM9Ei2aPT7zOe/mA7ttCZGXupPlEgHnszgyoLjE/HsEuxu2l4sMEtlssWf
eYs3f2BBT/ThW3k60DYwOqJfIUmm4NoUH6ph/J4Jt2GsfKolsOP6v1LKGHNsbXVu
sUZPwCXBEzSBxFSTidNhuCUyVJV57p6GU/nBy+I5gQGuqxqApFwR2kgg+aldFpbN
ifIq57a7VA88Ob2vT3cthmu9tkr2qj+fv4kBI2Hf90UgejvOBIFkAOx/WyTu0RYV
EEtD9OtDM3dItrxb5IovogZuId2dCG6ZDjIGkjuTwuwuf5fvKnzwOvioMRUQ3Rg3
f+dicIlO9Xe35etDfcNCNNsAygPvz6+HhsYwPyEXwBs2DluAqFdyShPyxln+SmWG
yVGsmpidKUB3LJJHn9kbAEN/Cwh0HWUbyVXg2IhUvrFf1L3tp5GPkK+unL/FLZf5
1jL1qPoSMg6I5STjwM+zYUKUNt5KC6XRNuNqXA2w1f43ocptjtUXuwCePP0JZMoj
NrX3uDX/TLoV+BcgeA/u0Ul1iXz8sYl0YxPhYb0SatLr25y4Lpfa/uKkX6rUkwvg
lXdFD0PqTG+4cUD2eV76/t+ShsXbXbjFtyfYsMOXxNgKOBQgiaYW7D07sevPjyK8
W9KAuLjxOVqb29bmoXpPrvZ1MfAzrLlkQFUdHOxMMv7ax6py3fGU37lpzXb2fucZ
UW3ebXl9DyQWRJxfCvGIOGY8tH4S1GJowiqaicnfAwVgvq1A0vEyoYLTJR935tmv
1NrDVDZvLlM9QLhzofvR2goRt1/OCEEajwSKp7NQVQV4cPkegSEknWwRzVK8xVAI
yQ7v73Ne/Amur35aD9Oe+3U2qzTAgbRqeGqbIHaNgFzPGJEb/J+PAVjzezNWmep8
hZXuVTCZmClVVFrmKkYiHDbR/WWhzx9lxQ07WRPTf2cNLTLh3G5YIqiJ/+Vqm62T
uqT/FotID+KxwwZ663/t/ebNEAoc/jMU/ecspr8C7mswF8oGGnnMRAFpNGi00g+J
JFSoxVICaQogRwpAjE9hmeJQ174+GyWPIfsK1FPHeOZaC4AST2DVF2eygySBwB6j
ul2GO8naMxmbOPPrYF1hBe/t0lkenAUftWmMxQHyhaNYIXjGA5F5ktQ6VM8YLE5b
+6PJl5+rxRz4xybBSmTpjJyfWX0aB6NBDuf+P9dNqTGxTfImZ61wGRkJlOAqcn+u
taTbf/67tijiT/L1XLObcm0Dg5+f3VuIoqD6uoYLrom79RhGtUsiy6rxQ6kcTh68
TWveGQSp3W3JGhgCnfiloqTfyzczcABgMqoNtmNGs+73UGUE1wS4R+JF2Aw/elLn
lZsOBaxvFqqrRbl9biT3ZvOgTdaVfQXNXYbLx5z3sWEoct+6bJa9Vyag/HjC8nev
EJvvyXKJ/wy7mKPxnaVQ0+TNln2C9NGKNY48PwGdlkpUEgVvWGAJz7lcwNMYXJXs
hktm2auG8EWutCXGKipct2Hqzi0nbwfVLCNxjY+A3ArqsSYCQrsGTQR6EKAttaG8
1F5b8QjBm8pLX9yYZiExgQlRhcilpmpkv21y5O5rGuKs3sb4D1ANPcvv2sRYbQeX
c+ybQHaU+hRjQZdj3Ul/U2YlZAeYR0nBSsUSQNeivuUyn5EMAi7Ebc94E4zZb/mz
5OAFwL4IUkE2FyyiNie2iSusaJKPrfvCtkivhQXmgoHx2UJb0jYn2vZhVx4dKS7O
ILvaOsAfgaiIohNIkR5kAi7VGJ/R7hrbuMDGXYvUdRSdehm4rnUKbZYMB/oJyQu8
74ucLR7L5rUp1mC3Yon2CediZKOGTtafSTtsebKO/7TnbAONfvCAvEAtsBiL9FUG
oaZ/DUGtv9cU9uBaYcGGpqrnH5+nGMtwQfKwMmsYK1wurSaJAzS07/SQm38iq1bD
q3ZOstkS5WJ0Bfn9x69wLVveABpCe50/Iq1N0Bi7bBw0eydd5mqXe+ivV7/FwkxP
YFUN9gxl/ejWeZC3c4pC4uER5RbBJZhVu7J2arZxHDO7eFjANmgVHQK9dppLqvSv
IzWCE7ecnghKs0l65Z6nINCQUR3qTdGZrY6wMZvwxiWHwEpPErBcASHCX9rSJ0kh
ihc4JCoIzaJn1Ops7WYLJH8y/XqQXmG5zEd6DUkq0qFZxSx6e06IdupCCyzncia3
UaUQ97XE8tUSHwo/U6EPwWdX8AfvkdtqjH4zlzy/TdtLyq4NCjC32VQQjMIvIYdJ
Bq1EkiDNtntUfVm9lizWJ1FGI8+j+jcfsPoTn+MEaJ560sU1XMmV6Utc9a05Hz86
8soWMcoKDWEKPPjmEcISOu1wqX97jVGNMUDsAtoXa9zaDp7sBcqHHqNmWk8HA6K2
Wns5F0xMWz/DdFro2TbXVaI+S79egYCDTxWxCegJD6oa+pDoBS3IqVuGlPyOaQ+T
UqOxPwzD/ZR+TnyLCiksBPOi4Onv14VwbkQff0KIGji+F87ThQJWjOckiTFUVrFY
90+Ikfz7ctjwhOftQuH5OrwEdvlMP0qc4tyuxHEL80tZRlw2RRH6MocU+Yb5F0r7
aPpLzZwfnAEFeTYVdUabjQN2B/wmIRWbvQ/CXOo3kl8w49Mhsoy17lX9b7IHPxst
A+XFud+eAGEve9Eks1QJkP+m56zVjxjSd2hshcHzq4uQlTvf8QbygYFzHM8hH4e8
jpZAdfxRZpqs3jZM0VwZ+e50CQsa14kVJ6WANjBrTYmHh3AP85j95DGqXO0LhRBG
Q/rORfNx3tstx/mhoTmL5JkGU33RSs59wlPwNj97oUcGlw0mSrwX/R9RCyQlWGS3
wWcl66VwQHPinahAG1eib5yQn5WhgByzPAQLI1vZmx2TjQr5ZvSkZAqm/CQjZ9Yh
q9cveBpOdLBUAZkNKwqGPuobbtbDi/yr50p8CuK2YAm/DRyAKaHghiOoNAKovRuc
AYz6Fi5/wzV4yQpgTOj1/mXiknS6cRIBEbW3ujpshp2q859ydG37SmPU77MUOL+i
eTazvmXeLZuGZXs75rROYHjVJ49Qz2HTN5RRTFNuGU43X+4i/20CgviWzMVBZu8C
mPeuOUtNWRg08hdsiV4l71lIyzFdOZe+MdxtXIPXF3K+ZDxlMXpHzdo20z1PCVUE
eP6lE51QX4Vc40i5CsYclf6aAB6XCghmVD3s6KxQKTm5BwWPOxcld69mflm1pbZA
2WH/pgljXqFnc4KoHd9gpbXdkzZiiFoIgkq/EQMFSv28hvhlrckigtO8TuxFXgcb
OLZbhs3NdHIPQ06cUi1c0d2Gus0o3S1dVnsIMDjTKIGITBIgUXw2khTkwwZFOa7e
ZOUxl+sN38FsLEp4i87sUrr4IcmlihVFvVB0owQsVJbTjiMXARQuwDPlNy2fpL5P
trvZusgSet7Pc8V4K8dGx/g/ype1b/Hg3Kxdr3wwWw/uKIvhTb/6mNc4Fkol71BH
tU+7sInPC1jn8f4byDBQ1MfHcvB4vvPu/Km2moOMv2O7aVqqlSqAh8y6aKsZ9bh/
OEAglPbu5/U+DLcgE2WWMB6L/bI3QCEvNEetp+86Q5ICchJo/zhBO9rTMkrYImKC
gXk4JGK8LPRvcX5sdDaQ1sub6WVsB2/csz4BMjUHLoRwPOB98r3ACxX5AMdeLy/B
v5ZN119vzedzxAFqYb9gq8JiQiixcde5u2cSgG+H0o5c0rRa5Qs6OPfbG1ktmUA7
bWG9m3/UjEVGY4o50OTR2tftToxX/laOpG6dyOASNeHSdb1EZn12NCI9M1E/dZAy
cJcowdvDxd3W8yk09tSjZHgjMm/9CzkXE7Q7W7evqrOs+Jrkoz7zUKHSsKIYew7U
mtK5NuKUFbEHT6cv0lHJt+0KZiRWn2MQQnzhVAvxCaL57vW1S9MK0canw3A/j1Ut
LgK3ANfnkEVOKT3l2ihRUKqW1oT8ANiS6aVfzykCP4tTB1lvM1vQhC/+PeSuIs3w
8mfL7yOjk3eFUrnxTdWndUzHRfBh0U5BkUnDToOmH1S12E8E4eUHHVGCTzEclFm/
GsYpa4KMP8zqk6kSYW8OKzBPsUT9GwWZsk3vHN8u7pY3jP4bOuuK4g4vk5YG3L+S
YRjj5iX7d9XrYylZ8eVnBE1ytxiVrmxxPcIbFtr1wGSGZIVJe0OdLh4ZHADKyqel
1RSEzJSxY+Nikcrf9ayaVsSndF9HLwzXI03zT1luWQJq+HzrMfn5oN7AjQEX1BgG
0iskBcXLbyCV/TR4R0GgEyvZgJddaeHspQpJRoMKr9M8nuwZbX5/0mCq1CtAG+ad
kKKMVmiSIjlv8EMOSihjL9J46iMLwXpbPJvJvSXyLTod5axb2inOnGvIm/hpbRVb
NgDeaMqO/KMKdhF+uwfctyFpfmtAGowmp1FZudzro1xJgVhcp25pV7kTxozvelXe
nDjYoRb6q+csrAFuOgg0EX9mYxVom7CEAR4A43tg6HhTkgB589soMPzuIRwW96yx
Ij7YzF2qwIb6e32kBHva8bbBoaBbxBL598IQOepLNJcZa6EVbFFIAi3clYWdHhZ5
c37+JPqtg4jJx9taqMG7jgXWPZ3wGtyJiKvNuDq8I9KK7BSVbOrwzAgFZL7pGRMV
tdFQk+nBJGJ+nmaCoI6gAipUGDiqsL/pCofH11M7LWkNNtBCKF9u4Wc+ZzR1PM3y
CULbHi21p/ZPWAliTSaQX/wk+3a/uWOH2nXmRjeyGvw0gOB+8WUy5uAQSJGSVrh3
wyUgPEruwfcUv7M8+nOApNMEZuIpKFi/3s8E1AQ1tAyo+ApMO9LtMOE48J4BpAp/
oKfBxZ39eucPCyHopSMb8/uKLmPNhDKmMObo2I7m2e2aC6FP4kJLhLJ36L1v5GG5
kyrf84XirmiCwGA64U5UZIVoLpJanPGyIjFwn9vzk5HbO3cL3/FirPkHLADuBHd7
vVAv170/I6gk5zdOFk63Chhg7DWQw7bUk4byqTjpLrOKE6A+OOSLBfKGEAt8S9Jc
R++GdNUQEXV6jEE/oTQ51pDnSd7utEBAk3EVkGk4x0NpGVNqUvUEtsP0m2mzzHci
WUQphJKcOhRHtvWU/gdUnoSckwemHbZuDyiJOR5QbSUI2liGH+gn7oDv2WP/GF6L
ucoyVkmALSNBz9mhh0eY2Dn0dW5AY4WuIlNu05wJYULT5TR28FkRteC1TUVbDyxT
Bav/AwelIKq/blw9iP54HS2/92EC8AmgxjlLWCw7lc8HqNphMhmACseYA/4sgM2S
KpqsDN0JXk1TkP/5zWjangInXkRzRFMa5AOKD0eU9MRxgE71wSW8kYdP21jmbreS
wZ4MMxuK2oRsGGEbB5S+nvEN8qf4c531FazaDtAWlSZ28/NMdao3OR0mwoKV6E/7
Vwwjw3CyqRx70MDxF5yGfu0jJ5ah2RaDKqfEzrIoxtTr1vrvhjI6ySO8ZZUnSZLU
tr/FylfXupug24ltJ5/kzBWpG0x4tuOumQZM9bKotH0tIyZmDs9LJ6gB+pun7Yte
QOc8eNk2ahzzjcVy6ox5JP/NYCkth4MDul3yZc8qjLJbpG4mMlAGxQhiwYZgLHkK
SaP9qmaqJmUWPKRvFT9D6RcNleNo7Wl7OlU4xFPB8w/2KP2zufWc5mRAyLLciAmV
6v8tFOgoz4NvF/vbQxjalh/N6wr96VLpdY7ktjtlD+i6pDZHHbITUXK5DHCSG8ew
yK9fS7irlnUmduose88Ng6DLVG2E0Au5iG8ZwNTxE8FipYwcQqotHyBIDzngkrlA
aqJhrP1BvBsPqRzvv1P49o7GxLJii3DZxfj0FFcjf9PPIaqM/PqkNrcxoA2MlorG
E2WPf59xzgPTOYFGy0pF8q+Jjkr0+fld3XaAXoClOKRlJtHBSDBQ96fyO4w+estY
XJlipPh8nVtk/CH831TNLPGCDEfNDwxRhwhwsel6MX2deoN2hohWpb17DA+htBsj
FvCB3/ildOz6zvRs/MTP9Fa1uMZm59NMxxEf8VH3NqVTBLxXtanZYKlMvnXF7T4x
B3dZOInLRmvmQ1pWeVoPlB6GgwwD5C4bCHR3djDpfJGTmfnQ8gPopkIDl44am8rO
6xkA3grcCws77Kpdn87q12SbrSxPLKZYJNlbHqMuJg6TDe2nM4+ahe/fXsbM1QUD
llD3CdW4rdXXwj+HUHsoTKuDABxrkvmefBXqa20D9v3yFMA7KawAhjYhu1fm6HmX
DIvj6HDDqsq7UI+szZfJgqyCWUz4DvpEPMAttIOpGspL63lS4Q1/396ayWvGTWax
74ZdIBdhdz64dj4eJ2f+uFrJOySvqflhHKm5xbsoY90dWEHmWPPP+9aUmEAfgOBY
yHfsjooDCN8u8e64eF7HyVKqdHajx8B7bkuTDDMqVKO/YYCxec7a/vJ7ZEuuFogJ
q7sHCdymp/F9YTBpOj2+Zp1C7s7lkUJPm4B2f2PQm0VAokDowIWOH4CDEPkzB1FO
derWXDHKD52KRrwAkPjW1Y8UMjt7RtVXaV8K5i3T6bw/0rMcXZSvQ3PqrLi5mNEm
4DWcmm+cE2yUDT8hNgSrcTTZ0SFKbTMAATJe5VWKmTaeENPQqjsYS8VdnBy4W3/e
3ilc/zR6W/cVpK2iBLdJacWi1AkVaGhqudEep7j//AQ0Up4kn5dFaMq9XLIdjWAJ
H8RSlo1IpVq08WQ1+5/mw9Rk/xh00WUtscCboYzdYcmiaXI2FtptChy1kHE0a1M+
MY0/3BBbz5xHEStkTUmPuKcYZhAlJ1mYoxsJ1natg+6KzN36pmmkyUigZb/jnUSt
FKuWyh+UiPQQJ4Z30f3dsjKTrgpD428qi410Mu+GlbWT7jw/FERiMrKyL1AHuRM6
tsdFd3fz41g1XPCMsHX20AqoUnslCL1xs9lYvKKaiSoixW5/OQrlg0vvFas8ILCT
lyYa04UQqj36xakChZscfMXAbVFLpdo7SjoqdM8uxxPGaE8p1b00h2XHG6/dl6nf
Cq5uWLOeR47ppWK32d7VvVmvaDBl7ywWmyXb99/Uaw5/SYybD0W1+mlmjO6AuP3a
tSn9yxvMUC//ekj3NUeZaOVVjVNPF+s/mUD9L0z9DVeL4f1e2KjKeLd5pIb1FMjh
mz4DqAFdFiiKAUsrz3MktysxDTFRAXYWTAz8iGqsV4gl78DP3RzILhrew9JmOhcD
X9sv37ghN9o6VLsnwHe3hLaNJX7Ocs0bK7VdB7XEL3z2JuoPRp1ch19TH4S8LoJM
LoWg3B4yooUEtbBSGzt4s6o4Ihb8eazB5GxV77SHVScxAi1XdOMbyjzEQIBURiNc
bhUgzQ6TY3vbpSWXrGxSi3VbmKpUqu8+m6oG9dqKFzDBKj+Mzyrd5zQY3FH4B8h4
Bv+XFc/K7GpxR31jtUDr+D6UtH+HeSfj8ASDOgNBWKnqWcU8jQINfsBuuJv7BEPJ
ScfPLtGujoGsr9zDXmY+yunN/0SuXlcBRiSPrkKrzoZap/Akgzsn2l1L2wEcdY7o
7C7Ex2zJ73SQyZLqEHD/T+GKBJT9do9b1J+g9wjj4qp+6FH3iLG9pw2BS7BQoNNi
rzttbijjK3qztCLkdwDBxaH7jrT40hbcklYQlSJ913XhSQcGM12pvhcItgMdRSqh
7WniU9nrgCO+dK31KD5XDxC/SEsndncPK+eIekx9iI362gDid/ioxCsSfpGLKaln
2bRuNS9pXLJIL801qPWZsPe+VbUKU/ogO4woh5wfHy9fkYXi5otz4JsqD3LuGp0G
jre21lP/+kYadD/z6n3rrGSfs4l/guxp37qfW/9VUmNZsYD5/1YqS3pFgoFFUClN
C5pQPcVb4VOuxfmD/cmTJkOySbLmw0X1KC69dpROvi97gDLHm4cIYK60LLb22Duc
5jEutDNnw9DbquMt94EztRl6cE2Z7HU/PiqrxwpXEFWAIndaPPB2KiCgx9uo3GwR
yRiI0rZsFG24SUJNTSJHDm3SlmDnxkjpFu/Oo8njGfPE8bSl2E2ybr83GHz7Xiwx
ceKZJ5oZ17J/epo60wSvd5jlo/HgPx6dYED71XTSD3PWpvLvfnu2HZcwdEUgaw9m
lPkgZS2KL1j/2H505NpQE7q1byNnawJe1crC0D3yHvjs9ZMKBbETAl1YJaoV7G8q
Ra27ne1Q0hSdN8xryUB/1clZNh13CqFC++efEflZKntoa4epNFrtC+mzedNs3/0W
AYJ92WWy20BPmgVPvbWQv3uvrOXmpGl0nfqbDch1kRLdklnfnBuhl6TqqcDfNHS+
UPM8rLwtRRYLPTreFELqnflzfJckNOY9T9J0XnlxjeAXvbUMytOKnHxeGCMXh0R2
99GN7GtzAj39a/8CXH1BVOL5kdY66C2tL0fA3i60a8Vc2Xum+Axi+h4D1x0bpTj3
5spjjUGhqXJl6JXCzaP+0xUvX0bQpaDm9eyRLC8OgI01O3ODM+hoFa0tGH47cWVt
UPET1NBzGHfDdE3u3Iyfe0XAI71ciz3R1c2QDfghNhvYHZKfmpztl/7O2ITTKDh/
6nGyISk4GTn71+U/9cPjvPIAXk081hU1LpRnP49PMPf/nGSlhjUVVbqcrI007cBc
pFnOvZq6vWNdZcLptni6Nb4BredEsYv0lwBM/8t/1XxkGkTmg7LQHs4mLqAafP9S
dU33S4g9vLa8rTo146HW+VwiUxDjATzrcadgUf7mwsgu38hy9+Jf2cPDjiXulTyN
inKpISi8ZvmMA0RwBkd11tl8RDfrRpLTt0+EvTUWKga9IxXmvoL7RyKIaoSAh5Ue
ioOBUIMMHAYKFUoOsWyqxssoAzRRgy45Ggpyq6wCoxqbQ6v76mLKLp+oXFjNESlA
qI86N9rN3TLIG9T+qybGcuzQmk62TOKVwb09is63QT4ZqMJ7ZnKr/4PqJaxK1AXG
ax8e2+8Fn/ZKzpV05rDrjUKz301Bc+rLUk4oTOniwAystvbse7OAWoYWBgP4asHN
MY/P0MfegxiPaRfUyUKpw1D/EmyxmQUGKF127kneTkl6v5LX4kb0EBpH0ikvEREy
SfCzqS7JRRWI1d6mdHRQzsbS3xJh4tdiVK3Acz6B51wyY+MBxWAK8UhGTOys2Q/o
R2s6dIWJSL7vJYT0pa+g7m3Jbf0Yt+Lz1epWhl2mL27u4bbzm3f7iMPVX40q7Vje
KVij8IKmGkUARRat5W1OvaXjXhtXUHHB5JUDndw4F/35Z1gqsfHvr2dFVHDyc4pU
GRPw8mUJiYaKMoScNzQXRNsbzc/+QU+qQRolECIsGD33y0uo5MGjPAofKqrWXC5D
h0JU/iiCvmXf5S2q6RMnsNqzhJ7vrk+2KvPlsHZmlpA+G807mS+N0/rfMJ3p3MEt
SJzZ02VmDVUqQwB3n7Ufm30bhjG+ArjUgIJJe4w6cJ1WOPyA89qbhREs0LIkjDI9
5LXQU9wjMZ0cUGTka4tetthBzONEpM/6NusXFr3bxmhJl7JZBoBb8QKZzcdEe2J2
iO8pCAqC/jsETG8j5hWPp3M94shbZSwK156mIEfLXD8PcZ7di0ds4fx8Y9xDGQ5h
TGZOF6hfF+UEUEwFCoq+Vcbu3JVY+GeOOe0nHE93mbokofHAxV07HN6qhbdou5Pl
8aKgaZ/bQ3c20Qb1+MBi5v+xStHIjQxzkk9B9iy9Xo5M06k6wQzduGopsHrD35qA
w2Y9W7aVM9i90OOf1ZKcAv4rh2Uyw5xXqh6C/7z0MioNAZRqxYPSD66MbI7G4ETk
bXcoR6H1iCmONc52BBuyVyJs+w3c2r/m8lHslupqiV1LcZCTUDIqHzHB9a8lSYxi
XR6FoueL1r1i+exkJuT+ouc6H8fV9ytN1t+dKS/SM3UVibTk9up2mLByRKONJmLi
pt6NluCV/RezxkdbrKCHJHcg6Jx0hFrvmRLIz4toNWqqxyDyx9y09DRx8NYOY6fM
rMTHqfSK0FWRBYqTISjL3DYb7W3qrRLZDe+s5MvfoA8K1/QWHJC5TTeSSbAyFYr/
P3acLofj2zksVYWmHFuCkDUEaQLZ+Ee6Ss1V5u9wjFn8/Esz5LQ5zbS+g1x7C5fT
ICrG9Rqzel/GgGkx9WeNNbNKIYqx32PlZY4q+DJZfRR2Xiuljnvwv+7ZTC3CYRpb
4Ge6GAxDIaV692eV+Uo3cUlaljMVwYK8p1AkWXus6qNxS69u+e3FG01MRTPIoa06
a8MzJLOZ7SqVoaA+5FRmazjzI65PvvQh3AZqCyRKo5isn+WHFDx34nmDt4hA6oW/
27CaX5Qpz2v05tPW83MtA4ljrc5bGprtzg9GyS1Zuid4AGi3PZPa2JWVWEmMFNaJ
x/QcvlP9E/wVBGz28Oi3pdqigzyRF6fG7KB5230uK49Y4BeNMQG+eKu0W2YxUg9U
ZFsmhqIOPot/R84Pj1iovahNilzbWpz9yNMbc+yKkRvAZta0gkBmxbQYR13g3Wne
/4dJpxTds0KJgw7DazGfjGViQ1/u4dKdrnET41EVftobXdTlJgvHzvJZNRQCTVoW
KQ/NF4PWETXVwL3UxlV5L+cq8oazqzH7j9IvO8kUhxISZGu2EiU7dn4kiQ9HRKFG
t1B3dNzSwEot25GQseNmFUtggnSfXRPpFS8Ob0mVGqlkQZZIsl8CPtJSdOS4653M
ybvIAzlyzMq3sIvxmZQPNKc6T/2cA8JQdOGGqZriYj0n1VL+rAiyVeHX13z3XZ+/
hiZZlvb+2jxqogSWmq048ae45BCURENFn9Yr7A3NCA6pSaI3spTmZvVpHqiYFmsk
+y1yhLwpASNg87LxmW9UQIPrDfBVbEOX3zwoQ1448x+cbjo/gNRmlK3+PFszexfH
ABZ4z7MMBucSN6oeQw3HKhM8vJge5hbm2l+F0OPsMrBbkzo/UW1LSF3WMfKNF8ao
AHn3ZQME+FoqLCkWonWlbtqONokMa2gtYnxJ4GX+mvTTI+YdJTvaK0hwBsqmQrS+
pPQjeL5jXkUzavhn24vH1MogO3ygt/9fbvZRGE05n+lOuYpDH3jbH/Z+XRhCw2iQ
2jDfJhsVmbIoQg8Zmula5/eltk3WzADR4xcbGkm7jYN9vQlOkEB8/x8XV2EldwpO
xgU5k5GJQfkiDhzGpV4V3A0aCK15kdnzzvYAJIXX+fg+nqbveCpD8Dh57EWbEBiT
l5aS5WkSwHVTaJpYB06he8sNoosHoRXP/JtSi16BtT4VO/DFpJJ4X5nCCnxtHwSc
/cqygDrqM8XtemD7jJL3ECcHwMAXxu6tU8CG5FvjpZbZBRe8ENTksKS7Ra0fLAr6
pGB50QiQBMI6Qp+3fp0fpp9qZFK5Butfc/VVEG0mgF9kkVDVU8eiRDzMCyh3YWty
YrzJwwfdHOs3XYD5CVCR1uE0QYq4kGSJJV+0FBAoeeE6pXANwYIlZRuJBlohRUfA
ahdP035LhFP+KVYkxhBZ0LZJoAWYcn9Uu/NK0Q7unkfihc26fL0OQhP7djhHVgS1
q/NBwFvPV6tNX7B3xDdXpakRhpyb0ulo1n9JXiz3Id2++ivb4N0HtDcs70rQaa9c
ZFZMPY7D1dfCrH1V8PPjoYhqhZCthmh4Jcn6RgSz3UalWJnjMFWGdyk6OVFX3UK7
wkHlWa1wiBGVePNFsxiqqssoY1ErV3aX4w6tV9EfWdyWsirLePz6p/pWX4abxi5R
+6vfPHOTRnoKiHxD1GUMG2/l7yLP9ggzMZYi5PYYgH/gLNfYVV8e1OZyvx65zX0o
2fBfIy8Tufa1y5ISOQOcf6dwpTB4x0genFzj8IwSA2X/xIkS2nYQdsJnu6XiP8qi
TOyk9xPAFezIcHGdfLHyg7NRNzfyIJKDsTCXQG3MzdXmRcJgWkaOCzfRPDaS5/np
v7w39rfCgpt4wXoTaxHrBf1C/o9ZO/pe83iOsk8BMcO865yqnGOBe08f18AP8Vyk
cYjIye8IkzwaePtxZyod+b1sSmBvXvwML9QCm9wZOLm5J01pfPtKa80XJ49n1lhX
2JFvehG0PS80C5sdXeUPml92S1X6cPUTOrs8TZ88Hm1wo8SffjE/oGizv5enalRq
yXACR2ISgnd2jKS/yMfFA6f/uzcxDxFKdkbs7WTUBifVrWw43OlLGqq//hYAWhOA
WaL8trUmgBBeEFUHkSce5LB4Fe57UyoHO/eCVwpIWXl6eACVTquBNUrLRMe/SX97
Fwn5NIGU/yos5CAKbPA+pEb0hYxg3AoEZIS8lQrr2cd2nZqwJcTFF67iNos+QZpl
MGZf13eNBL7d2/L5yuoFyLv80DmqNO/NRaCcSUOX45npynKrvsVxuA1gGOMNDLOV
Q+fiEsgeRb3JU42FM+S8ng00yrpMnxu/0tJe6b6Yh75B+CaBupgBiqFtwGOz94H4
pfugWkFjZBDSwyV7moq8q4PiKEEXHssbUg0pJRT9f1n07576XObFtu+lPm/t3+wJ
ENkWQwrYX7+d7Vb68qqI+t98k9opbsXFvrcAstLrYRBCKo4bLhv+yVmcUl+13HlM
Bp2DHQm4xI30sExEhGuMnIqYV4vaN9tqvK6FNwt/MKYGuBAyNpoIH5P0KCc75pUJ
TQhEjX06wRRt8pdgT/P+Z9dA2liBTSoIaXayGeQ6jIkW5XBh9vvq2/fSUYmohaTz
ie6aH3daW23ilfRpKFYsENtXBKRMiRLfv2hBr/5jhXPE/kIWYyfYkNRq3rWmI7hg
823IELmlzhFcCmKDJFOweb0rIFvh+gsNWp0Hbjhkrfz4aLKht0J7MCUXIxgR6Mgv
qlZu4+49MrrNL0XNNAwoPOWFqG7Jigr64EvuIp0jQVyhjC77xDl5kSBR5g8qefp5
uvzNyoH08gGPOUohGPIQFr8JrCm4mauvlfr0UJMj01w4Q74OD/i4ai2S5gH4M83j
mlCR39fGCPuxD0tCsoN4AY9iQz6vxnwkDqFJgl16xzPoy2er+Q1N5IZ5HUwDQcMF
vi+DVfL8aufLvAz+NaA+N/5GFnNVdexy9453ToYvP7v177BbPe++kjkreiH6xxZQ
Kgw+MnFG3nTElkeYoC2jncOSUjpCC6UF3E0c+ZxhY/tIUJM7Xz7vZU0TNgaiKX9d
Ehqh9fnAO8vwfjPwnUhNQpMcsZYgr3bw7HS3f0F4kpEuoM9yIp59CH2l4SFAjNHd
v4k6AUg0gCpkouU7wy4QquB2fi7/grYiTxED0GrxPVYDU+OWPQIU7Fb9/q7Xb3WO
tThSYEsYhPJBY213cG8MCzP5mjHIR8vUjDssuiLB0E0nSokmp9tDj0bXm+ogpQwr
balorYz8bvEjpDJCiE+AAq1E8JJQUBNlyf0s45IGIFh4EFJUSRz3qTBiV2GzjKDH
D5UGolkjYuQnPd3clUgJjw==
`pragma protect end_protected
