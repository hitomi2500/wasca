// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:20 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qKiY4tWrOjsOIJw9sPF52R3sD5UuKFndpSv7MIocFI8FZaNwksO54pZl21L9unTn
rDf1TGzQEOsOhay0+dznX7vaUy5+IDlzr81IzAEOIXY9Vy29a2LTY/DB9VbWa1ro
nWxzSLAyuuwDen7GPZv9Jtxel9utPcongL4RMPWTEfc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11712)
WREVTGyxpEhIkcZR6BAeZrjJEi7sx4JKB6H5lUfn2CxF2reC7tgR7Eb2i3Wwvo6x
q7nf+tVmqGKXp9FQNXOtVNZQn18/tuffITfLGT7OfmRNTn3DL1S+D4J5yAVOC3mo
PeGbO6KGbgSusjYBoCwRZ2yyRGRhnKjdgkwv0I2T3Db0YnmGltXW5DUZ7xg7dd5z
45qlAFkYZ7ReK0l88vB81F0xLOoodG+HVv4/OK8bJuCAiXijscmqwtz1B+9tnV70
zMYj0B2cpw2+TqS5bRYUIH+uvUzGjCIchWRefpR83zhywS8rgxsKOrk86puSXwxI
352YHicDSYe97N0URhyhSkW+09nrwPVkgkt4tdOgxZxFbKHc+JBt1S4VKhNYLUR/
4hx6optCa4yLJoBuyRWkqjtBsVM7bamRBXQEeHp7pJDiUG4etdBJEt02b3tQln4H
7H2oHSyU9Oft6nVQOHkUCOgwdXt++MeRh06ROmTxX5W7ie/+RlasU805irzvUw7n
v7cV2uZumza/kW7mVOXiLnl9+3VO4azRyFjxkE6SoTXL5JyiNgnWlilNKaJd5uC7
LsVUhLsABj/iXbzewmpKOF6qan8bkqe9tWc3e09mu/rNVNP1H20JmmblGAB0GD1c
kUarwNVt7EPW21WFEWtkaB1ImM+LhgOZwxBkHsbBPv4WCI2lN6cidgsROz5+ad6u
+Rv5PJyhB0Xh6+gmpdKy7KpIJyfgRG57CqxVbqlSK0jhmsUpOp1ZrAnXJfKZBDkw
H5/tA5M7IqcDPE5/cQdspTv6Z9v3fQBQKUjpv/C/U7+d1n3dOMJfkX+9A0yPOtrW
HnHfIBLvqmkqaz+dZfAG2ooMOrnh4gQlGynD9M3ANGrWVBpVyy7+RO4286AHVtjA
TffsPc4vnxpVXjNiJv6e5S9dvszWtF/bSyAtTzZ4B7sxfBexu0TArDPeGhLs7Sov
0KAQvJ8FW5lwyKxVHXqXxQFEzakhxSUJGSRMbMJz/FqCbCJTpMN5Rf2bNE442sBX
MT99G78bAzs9w7xUlpb8hqyz57dlXtmUsc7/v7TBF075d8OoHiDx/bH3pd0S65t5
rTqRkzpqwA0hR7EsOfitWLRcYBAH2HsrKYdpaSaT3Z/qPC7EpW6NMy3F4EZyDIJv
+sbmBTZ4GLB422JqiQlVaTVY3YcZkJHcbgSJ8+DSUgPq/JEAT6+YBtY/tJXFF55F
d9Akz/9xYE6z2x3nFYnHGGEPzRJjQ/Pv55DqbyF9sXqFQP4Rg3YzJhNCedP4geiL
c//i0KxR9Ni7sGWDvIF16oUhEJL1ZqkOuGTHvbGV243d2xc1NtFXJtYzV7mgK15m
q324z1MNxwLTOlaw7GUO+AUhrKP/ZTQ6So38fgIt4vKmZWVd4xOPiBZ5QxprmCvr
OPpX7vOcunq/eidtFq9mF5otzeWeiFb5OzN9kLfYl02LgwUA3nuFtjJFomsS/MkF
hYLWZ+lUNzRBGPsFVHgtFaSICsJxpnwnynvR1LprZZRMMowz3Y3LdSHgFLHjc92s
58Bs/+1oNP9G4Q5l5cHFlppbZgphbmswxBgIoMsXffFlLKd9ayq+L8rSbzZlbgNX
MBZPn3cQ6T8diO1EgKPs3lPDLJ4i/xrFu7eyjl+60OtFc+/hvq9Ob+HIn/8x/W56
mQEhLYm/2pIXAgQnOTh6ftzBcvIQzvgAHaVpaAANP9lefZFd0wmRi2wo0R87aNqb
QMXMke1/OAi80oo49354lHK0BWEDcUBzdnfcAepl+yG/rPYRpR95EWIFrhfVeUaY
mW1ZFCj/8wEnobL4TA/Qbwe9aDYucnl4ssEin0jzGnzS5rHdv9zm1EgdzqkmlEFE
K6IFjThCbVhR+97jDVy5Kh5W+3nmETKUUE6vuicR+UP5R0MW/W7Z8s3aSmoH2gOl
FXVtxMWFH9deqy1m2S8J2JSkQogUUtJ7XGY3t319wHqKJ7ghp53KXB042BlnHvVl
yp51sGNZHyhI51I/evdgHK61mkXDOaPUEhzfFJV/8/pH+Xl1ErEOBp+Ayhs7ksmR
w4+6vN/wgVdsqquZJm5uaeZ3FOWfXj5GClZLWTPSUdwtxHiC1K4HL3XNiNUoWZ78
/QCqEuAP1IBhDbSkEoZlbkFePHX/jCreiwEtS8fWVCvjXf05P5Pm2ldZl9Vo5/PV
VZ13jLmMX3BtDXtW97eNBAyKX/UDrlYhRsia7Uc+zKRi6VIkGvbvcSIDDt+v074n
wVs6V/XsIasyGd8OnmydZe6BB97r9LFfGVq/obbtAIuCEWaia6f5sn96q6OOLH9M
Z3zPciTuUK1JnDVwRatouAAo/0nPAJqtX2YkXJiRifEfOijQjVKUA6lEdhpp0NyJ
BjBs2xUZsRhX/sraM+wfqfm4JJxnxq/3f0BCgwNj9JBbauUrfE1HEvAW9quSUJDv
d+8TYce7CRMtZh/w7/3+b5ycFMihNOWe4Le67/j0Xv1fKBolS+ez2LDNpMqr3Am+
8y98Pmzo9gAkvXckx03rBiER+WssRMQQyY8id6CjcWxzgL2+D/TxJ6s5yfdNq1C1
XVrL7EYKWHksWTSPyqrAScOFzAw4uQ18RxBVpafbmM/5TqwhcsJxnga/Y/UQxLaf
XB3w6nE5v5B+IzNHvEtBC1CAAj5go05gmlr85vtY9q7+hU3jimd3dpmPaaVaWN4A
wfwKGZcaLk7A9nOZY6eBJrtG5S1/9Hwx7C/yFo4iAzbcRxA86SWq6vQxLQSnDFIw
XAtD2SfKpLLqzFW0YhPT4F+tO1rxTyWW7Vv8YzPds8nwYhcqg9thNCvVq9xREy/z
FheKnCuQQ1jSa/3lJb2SgDvv8gMQTtT73JaORU1pbpq7q9/QWNW4lQ42O6IdIpaA
Q+xusx1GNQQISyzL9yAg7NNPka5knLsAaUlobpjSB26dMZbo5aqgK6QpCNKgy/9l
JsZDMzQNZ2sQH8jlK0Ax9cWRmCcKEigslLGaflgd7obwuu646c2jixUhDhLT7yiG
/Qx5+TSfWPdiNz9myUKi2BCuMxAo6cI/P5/0deZW8+4FTaG/aGIILTC1co7eV6Ph
G7vERk6TicZTvnlQUj/mGgLDoV+ZCCpjvsopRD129X51xh701RgiZOEivfYxHdFF
/mMxj5pm3j1F50hM5l0FM8ivpdD7LiEaXZzZsjnnD9QHDvIYVo2STh8yHjB+0I0S
i6pB0VnkDq+GKiLjUMisbRN6640VYKiZlwDXAEfFJcU/6N4PArQDGp0+BSWbbkP/
AdH1DE7Xeb0oAt+pGS32REEC9JOlhjOS7q/UYGSyacfuOl1rgtvswvqH6QL4dTnF
fX+POBakUDI9Qi6SDsFWwChw+u/MEIQKZuYngDRM61XaHPmBsvHzS5nIqCHgzS6k
aXUZddi4xNXBCS/CMzrnDEfNrZEBsX6gwpUjuPtshKhZRjKf+nkohtcW0UHhuwU9
MZuy455M/2q+80AM50UQrKJ8zM/R9a6GHcPYyt/TDGji3V9WA5NaxGIyUJYExeV4
DOUrEBFVUKtWBXlM57PgEhZbxrNDaUljrpV+Hq68bBIZfoDBlW59tZExvY251vY4
OrlJTtebKGAwNwhfikN6WXaLeyfbbgsWLPu57E5C4uYhmz6YvNSt3eLOLqnLWAQG
YzxrosDs3Gyx7liTWHZbRYOqjf5sn7N4c2efejo5D2eibZ+te/kALFVTwbgJiT4s
T5DmNBu3+VmNxiJ5DhVVDq+GQwmiq4UZ6doUJzmobZ11Rg3MB5JkvHjx3oBa1S26
d5K3KcJqU4TiX7rJ87lBw8FZUJ6VaU/vKIjLYX52F9v0VFH8KLdu06LgWxrc8576
01QDZ4HEcctBO/xYf4G0krwNT8Xe1zz8o9hS462IgQ2XzSJkDFY05syHakkuI+gB
186tgpfc1Ea0xkmSxPTelhvlyLlbqDRYwmIDFnZx+TsMyPdDrkBz0xvVNwA/cP6O
pS6l33/ZowOQ941AtnBi9HGjP/9hf5Zd4HOhDhkXxzthd9qGioeDxCKcqHJ8GVZo
3trTJn0XxgGWBiNlWY9355hJjnLu1EO45tEZdEHU22gQpL8bPwHJluYjA7IH+bRU
YdbbXUl6g7I/MqHpyXRY1jOxZZcRADZOcuYLwtjTtIM7Gcw6n9LakFUesMcLsvqs
jKPGCFhZwjJCT2YhwaKzcPTAJ1w0wGf5Y386TrVXpxaKfpuqkTWxw7EvYoCZXJIL
NPIeHxzHdLFCqDG/zuwp0nnKv8XgbWad0W2UmacgdYw8D3lktt8SsXt0tLJ/0FeF
gyzsEk8RPyjsuIE8hVAEWBq6gb2hS3NlOld1up7gDarFRwAxE2Vgh65+j7OcLvJ2
d2ROZS++Jsn7CNt4QcyJhkJDVSwAC/bHjP3jDQvZ8LVnYs0Wm9cNASJjrOPIyA8M
fpNpYGkTzCiWmwvqv9+BBEZR+YjA3+aq5I5+Kmn1SIREx1k1+ge1mtTNYN32GE75
pKJpvI4Qia7EhdYqFJmIN9lxVmx51SzFop3qTCAZMQunY/mzmhM8buRl5tI5gb6H
qDZbalfMe29lo0xDB8uFmX5pJsPnFoS2p/ro/rzQvNYxfdU3cFedb0ti8wZoq9+K
h/FLBbUl24K48NNkkOT2NuVyWb26aLHT/7H4dLCkOVWVimFC7r+P6WjsIRNVUkrZ
aaRwWVNqZJAVcqOtopPp5jRh8zsFbrglRuavbCaRKZqr3VTj5SEMWGpAkd8mvhR+
yVV6s0b3qFZeD/SCsQrvP4EVUekz4bjw8Mx+ULtodSHx/B8eTzbdZLhU1lxR6IwQ
rr7oNeXqX0d9dHP2aBY1swZPpbnjLbw10gQZIFoW2NLLqXoma1JG24fofEacqSd4
ATLbesTWmOjVX11J67eKDXFMRGKskfAm47bqxBypuBKBmklpxXe6fQvCb/BRq2ho
RrQhZW/Y08cCpyuuibZT4AzEKuO0OWSNKBlZITDfgYi0RVjeB2Utvp/bTvmWYjsd
49vLU8hMbDQNzbVjjwqbVXsk42T4Nl7NNMcDUclVeiWHlZIZr5saEicNtiyPE+yq
j0fgnZ00Zxd3QTu+BEFgqmCscZPK3hLpKJ/d5jH/brLE86UxOpYOTg8aoGgtBaHE
aIxGHdjAEzD6iC/E3o2KuGcw3IcxF/JAvNZZmK9Wj0q7W5zBgNoctZTinxH12wXr
6+sFIMnaEQD0jcM2pcWH4TuKFVEItbrD/r5lzW0yEYEuXC6P0DlmvODd6uz2TIgq
AcipBxctclMvHR7H0Da3+0hF/NAwoki46C8jUpiyVvY/2iUa2J43Gnqd2q7dCz6O
DvjQqDqQzlubSnz3D+s0atohxIzghIxqrXhzB/HMvHF6G/MWn18mghhwDQ5QEJDN
QTcRQR7RjizvyIF9l8VEMa50SgnJO5oaWPDgaJzcbCF6WlzD0J98Qn5zPrMM+E56
d8SDmZZ7bIBDEEgfO0m/7pqSKzmU4RfAeXhnLtCSbtiCKbRmdmmzYgbz2xPNf+y9
NESyb9bNKfvLw2icyj0yJIe5qa3D0k4C9kBl/I1isRHVOa3Nds6SfzkA36DMdikn
5QQ+SjpRlRi/Y+bGOk6Go+Dy3ZKXFgyrcQGuWNKAU6j1uK/YfgRIKNEbnSz1gDki
0q8XyzyWB+rPBFztBev1JvfYW/iWWOD1UG+60PgnmIfJfxO7BwCk8zvbzdlH7bQO
aLTH2Q106Dt4KdQP18w7lOKogv2AwhQYgprH5N0KeTiQ75UVdztmHpKDOmPjA3EV
nXYLnWybe+GjsDNT88x572MBH3OpR6GRlwAKxueh/jShKbK0KKzh3nfMtLhwLKin
dsWH5a8on3z7FlW1t6KBhYfYdUc1bt4faLqwRDuiiPY2dZnhK7DsVqvQmqrP+NIo
zKV+PzotHl2nOIt/WD+Xa/W4nw2AT8kv/eOrUhQOKy4mRImlw9HRnagkRQ5dXvgR
1rJoHYrnx7MbXNmgrFxHxDaZfty8/CFn1mLZPB3HdvCS36O7RORyH4WHoMKd0q4n
iiFSosD2Ms/hBkTiOAu0+zEO2hAh8oemyoQlxkeOd6k4lUB4bP9XpHJGuUjOr5ro
46Cc9feMbqB5BNEADArOdzCh7/xJXcxFyuPunNVGHxZpc2OI8F5YEMqt5vRa2Ttp
qoh+kNLpe33oeJIyESspn8dkqfK6vHLfXSeZF+Tm8IknujKYcSp5Y1ZkaDQ+e57o
7Pkx43SzZENwpQtlTz/zQwD8i9RwQkzrcMI9X4g85X2ro7vkC0O+hFjLs5jaM9Rx
Fr5BImuiP2GbeaBSTxkZMRPcuEBYgxYPweh8T+7OJRlLRFqSwy8dJZfhtC8r0QPB
FrzL+HtK0QgeZO7h2BTC3lokysHrVIUyGjfldb9vdtlGwzH7fnVYAhCNJhMqtHy3
j2nuulDmxODy1L7drL8j3IJ1sl03T18FhPZTZHM3AO5uVKYpI7UGXPJ/VFtzv5ly
/mw24UYkHEASgLm7HPKsovTjVJavnUrj1XgdeFFSrz91evtydUT87gXJ70nGk+hc
AkG+UM1T8EoAb/gYy7QDQTExJnwY85v2/cbOVjcZiBBBVbKryXum1UA4WkBHniKW
9v6/9oskzAsVjESAIGOh8ZiFmusooB3CmNl1OD8O8RW/aX7fZXeANXVn82CYlDL0
pqm4Ac4DPfAFDPvlFxiS1tsxQvBYw77mTQoMrJxUN2umjQq1I3XthkVGx5fLEOVY
rXAe1m8u3gy+cKXWn4Yii6ffgW02L2JSkGOTh4BnrjXwhe8KiI2kDpP0LiNTE/qi
dJjIRapwIEwAWlzJA65w5tDPE7Y1LIha3aip9nKHlVAxXhK07KBD5Kb7Do4HGvNU
UcN6WDP+DpGG8ePTnt8Ay8tYkLY1TegCGZtsbRnCZHsMxTrCtUlYxLzq3IkMtCI9
s6JyP7OKXb1/0xETwLbCYV4vEPt5zgm07a8q2WqHNSp/WMlsQC21AeEZ3lJE3azb
nIA4Rda0SlLQMzzrOh2BFSwYnsEvW/OFsSYpUhWMkDUdvQnZ6Uv7o4xTWg99TstU
CoyAjj2Hq51psvud0HuWg/4WXOV7Uf8DKv5DaGuly4oOe6D4faT+GsaCdA60Bfvm
4PpptpYCdYgLico9lTk1xPN6z5ISX6HxIMBmYSqXSaXV6vDrXna4F/cHRkF8F6+l
GegAFoHU5wwqKDg5OGGkuSL2X8Z3puVEeVctm8jzlaMJvZqPaFdL0MOh9jK6oTZB
lD2xG2PDWBVLoFgWR6xCmMwE9QBxACVO92LQrsuApWdF8+4IFOvMI3Lq6ciZ5xhA
FDbQ4HoucDvnQydBKq9I2RHGK7J8sq3WnB9WYQCeTmOJBLN20Mkc2bgb07YKgpPy
UjkSEsHQInK7v5wEqIOJTB5t/tJeDxzjrdCSTdqsPr/fCvHnRfpHFT4aiC/6JMKM
84mLomYOMNGl9huhtlRnAE9XPfJukKS+RVNu3jIlg7eJUbZe3DF/mS66amCh5YjF
eH9havRILVc6MXuGOX/TH668njrIszUL2WL+e5dkKNMdD5IVEdYJ2WnStkgoP5z/
NdqkUBf8ffsBOqrN8CLAhvV4G02jkO4F/XjybGr0xfljUw22OZgjCuzLyQ9CJFr2
9DpxNAXIua0MNLyupcr+O0ZsCJ+KQGGg/xk7ExUjYRgF/zT8fOaFyUti4hmdsGdu
qBap4iJSvXBMZtphjAFmtDgsOuMWsoLgx3hytBEKbrUOWWljXTNJPBOQKdKkmT5l
+c2Hm4ntJCMrCFYiPX3VRlsGkyEEutHmgCNrk8svtYjinhBDjqQ9OsnLXZmkcyfy
Gwqckfhd62hoaWMODf6ejPyO1dq/rcJJGtMOBmajtBC6TxHjvMBqYRDAXI/ReTbA
tVJhyH9Yk1FzB6FNcIr5v+uG+pOsPQcIx1BlzjWQYA85hCvPbYXpHTfnFJKt3oes
ZXu/l5ZnUUglhjv8AKthSkn9jbgVjDmvzdE5/gecFbqeZnbGaTx8pgIA/8vIOFoL
ScpweyZxgbYZtHu2v4ODbVBUiXt2AT8Rb+uRZeKuIdDCBSpr2HbXcgauJysNjhKk
IsWsYhu5zssFjqr2ZsW/VGjLzseYAYF9ycmsqKzU+5MeZahCu8VAKeabg+VUYy/N
pmEV2j0a/r8wA//VpRY8BQgCMUkxim89PnnFGaKlr2i8+0GhhcXRfBW3xArPWp60
SV0v6F2CqmcpgYveLZsz7q0RxmAGzQadcHfNUecq5RRdPb0/BqRI17G0W3LjjgIq
y7NMfpf4fhn5+/dS/RaYiY3/HxvQv8kaSvPSPw6e17rJnEQOt27H2hCrhkHyYpCF
V2D12tP7ZWDbszRlFIxwgRj5j43PvKjURSQ3Q+nkObXElyLaG4pINw3tED++XC3b
ok1Iz1B2qWYr/5DP1yv2xgOUiZUQRBMmPzljr9bcf/ciQ9Wmg+vihQunHg9rcxuA
eSpdu3CyL8yizSu1hfWkJ07MO+S+K2YNzDqvZgWS0ZHrATnbR5wkftZixJJ6dOFl
afdrFG08ePIfN5w9iu3f+zAdTlzTzjOJMXFGlKi7kQ5vHnL8cKqfx1LIFBz0P2JO
ZY7D+6GgpAmuweewyU/ke6pP65jzbl9L44EIM3JN9StHTSk9uGeeLjyVf5uivaPe
Nrda43mLljC8j4/X3BDGc/u1gAsMqNGi8maeTg1c1BUdyfy1i5EliCKY5JdsMxH2
OLwfHn7DPNkujQdm5MCU/pkjxg1bn/k1yCQqdMM6xHG03AkHrg9LPRD92lnLWNEG
0qVoahrC9qoDNhcoG4iJZwCI4fApSb6cyskJ6FEs6YyIhPazNuHPQ0AKYlgb80Mu
nhEu6n9iXVmmLfg3LeGVWUdJPp0YcAQxX9lXMOpG8Hlct3NMU9QcAwYCYO4mWgXT
rJD0UjSfcHv9fP2fG6vgi75MIXLSwsNmTi3vdqRGrTL2o08JnRHORVMOyayOnWhR
931DRKc9uDnV7QrfnahZq+ptsnmIpbqY+UhrF5TzneULPVJG5Kv6w5ez+o4JoOj0
vOlJw90A5Or7vOENraNqbsSSWdxemxdusdSQZ6DmAOW6wMy/yDdJi3WQuGk7uXLg
s5EB8HJR3As60kYIgEElvThXT46S6PDjh41Vk1ww4rgwctpCubjp46SDi2w6Na1l
3cYtJP7NudHy4QqarUZn1/6o4SiQUtBla/ugbGAv4DSZl0IQn816LIeLypGQxwro
lqH+LJwzgajgL8Iu7PVvYZs2unbO2kkB5zCcR28dsoJoHZZe/wEc6sTYn/FyDsbI
1d7fYJCTOw7QrhlJcjLr3z+J6cWQtEqNy+bEyok+4YaoMe1NOGHoowpx9m6x6jH+
X+NwMnlMo7y7X+P7ZtrLDHgvM2D8OCSRvJpcvN0RVrZlXWUHWUkXZQkbjRm40pUl
wYtqEXPO1bvc3VX4jpupJUxfAgZZXL4ZNq16SGUX73rKoKmF1C3RO7wHNcwN35AF
H3yIxa+WaRZLx59hZRJmVZbQn7bEEQatb3KZLJ5mx0rk4n/c9EakpQVUMP2c7avz
pTMrDcKaUqXX22mMcphjWWE3NEUnhnGkF1BTW87bNCV8cZVLQqT5aJIywLneOFnj
vURaMdRrnWAjCKHrwKHuUWtnHf4dSRB1PtDuTqxv3F9eZbbMzS6f3IZheInAPAli
OwAw5E9bUYyPgFsPl8Q+8pWZyGkw3gjJDSOue141lGvCmJYRinvHOvegVfM2ljL5
Cr2JoDxjS3wS4MB0lNEoDChEOjf6VReQ0ls9A6cGgUbstxV2UeSMIXkEJkcBcOnS
o8fyfa6/br5U8jqQ5zOuvwAKUgYDNHwHzdyhHCDhzB0HCZzF7hQDRA/R7mQaWRa/
lPlMpNRee4GCKNsZ3Crf/xnP5rnJt5ZN99stbRa1AJT3pJDXzXIk2RINtuN3gG8e
4YzegXx+VWfx9eBx+QPT1vVWPuwG7a+BFwOzBA7de4RFZWQwfZsV7jj2rqBK4a3e
mm1fBt8m1flanB/y9yquU/krsajEDcr6nG4NnvfjbxwE2iERYinYqG4E5PZ2jkoQ
wVti96UOoxlyxqQEFUIXt7kB8F289asp7w7VzMUFbNnVF+fFONCTzdOiUtuuIuqb
P3uFPwTEphY869rcmlR/HFm3vebUGsowPf17pbc7eY9PYfq7yR5ksef2rn05cnJ3
iEy0JH+a1XmkJiVV+KcwcmF53Umy9EZaYcMt+hpiD68/LFDJFDCQ8vaU8qJJH9cG
9dRBUP92qLs9//Bo1HhIDpg/ffvknZ4888qdPdHTD4rnjRitTPhi3dFQRTHZeQ0T
onn5tJl0FS/nHIpphEJjEtWfJzLhmbRVJaZ1ENz477dt8u5MB9rM+EKxjP44uOFy
zCwFyTd16FKvhEc29jCc8AZkNpgOHM4btB2Xj5xBKq5/2MBz22/8z9/2ZshaTqPM
Hpv9U+MtJlJWS9vGNordMTJ2maZoMVPqXe+boF9y0Yy/FK9ldI76IalmSoH8Z5+0
b35uhCzLAl5cJAAyu05EUC8in4u2s9b+y8UVYs/AanMJXulRVaEAqJQgQIMfZCWR
nHSwpBryDHTz0owKsIql5vjaEkJ2bubb6dVmsiYjuDldYH26NRYArxkrgW1PFRUr
MuMgei4xRke1DD2ZsEzAMAbeQfnHWwHzY5TyyhJGsMNzO60MnYWnNgHnpmebVs9C
m84OWeCgbAmoUTTP6Fwwr4R/q1x0USNDjes+GrPKkUQ0ApIG4m8qUoBQb+e2XcmL
FlKyTReDwfN4FZi9oLAFr2JUONIs+p5kfiE90qFSzbdYxJjM37+QHxOczu6+4iOj
EIGZIMctiPYRlYzT5Ip/HCPdOnC9AeUVCYsnG+EVdECPu2mCL8ptabHMYGXqFHhj
nfcfuN4U/x0QdJaoSwRVlOyZ0OuJadfDSnJWxrTscxI1cTbCiEYfAgKcbFIJ61JT
VZwQM/iEmh4zUq+E/fboOoLeX9zCyR1FVwkXZ4n0hglM0fn1HHyTVBi3PODV7jOt
ySfUPcYnsnQFqzbZYslcek1af3ApsqkMUrxnc8EW0qei+QOGXsYQM6af4RRy6CIM
kyixomICAM12llnnpsaxfFpyhBYhbQY+0GMhZ6L6mWdpKRRpynK86rcMvnxLbNwt
FWHJwAfBpg8iJsmEhTmnTUM8OBRVR5nla9N4+LpRpQ4Lx+hq99kGDnzxrs/bJspR
KzsqINpwlm6aqth6ZRXTm20TJz3VVaYwtmyuwTOngokTKDtcUfQhW7+nllY7tUF6
2kQsvc8wi7fBLT0ZXb+/r8Zag6FtO0WeL/KHiV2ys53KXgiK0jW74gXUzfMjZWIx
7L76jtk6wAJsy1bCP9pAHN6mnfo5CAj7wb2ILzxslQ/NYyIZ+SuBxbqkODo3fxSH
OIRKcYhh54umbTrg2t2rcjf0XvSgy+Dr+au4twIDuwLEhA/hYWxPsq5vJ5O1vo8J
K9vSDFe5v35GQM2MGY4IVhiRAWvskrs7tysx3aY/eLhZ9ab6vldh1MzWv57Nkbfx
sf5iveBuSvyY30AOjbFj9nfx+s4SDFr/sofQCM9z6utG+DLLPrz7RAmF9Mmtvngn
jAVZ6lvliGMyZoZ1U0vQtzneADC10HDhqYrwocjG/FWDUM/6HqB1s75BOq1ypasd
5+CAy2Eq/4ZrQWz7MvsQ90Oblv9f36/yPb4/ue8R/X8VFyPXl2MUJ/pRFt8mv4Fu
Srp/IpiAX23EYYGTnzBuRMzOEluAzAcvJvzBpx+TncalSH8+pnRQot77KPlNvBKs
RC0sX0qKd6U2Vhn4ewQJRLWkQj7AGTRjK9SkEkX9P2ZX3atme4AajWajY8TNGfBv
1uGWHaXiabmToQKclFOGk4R9Rb1hbhaEeUQRCPf+3an907jdPyHUUUNlF5uyE4Qi
iAckPIKtAJ/VXnHr66bhTBrejrsYQwL7ejV5L+XjgX7U8jip75kWhBWyAp3fCC7l
0DiaoCOCdByxdz463ro0L9TWP1K7HjQkYaQEAQpbauuOObuDQ5cMLAkpdDmLPBTH
00nNZOJ5N8oavR1kFHlwZqDxhNTWt0ScvnW9co4/ReGMA+nv3BA1QWdjd/XaqSF1
TDtdmBQvftFb6ndGQ1oKs1/ljQFaSOK0QJ6VEFsOqV6WzEhkobBfeuRN/zPvv745
FsVdta9IuI9GzIW+vBC4wKeNBxejekTopkhOTnSSA9Tc6a6ffMBj/2HimmOvQMcm
hZvvD2mItJrYzQVcFkFdvXryQScTl1P1TReXOOb9HeiQ0dYvf7Oa0W3bCpNFXxIl
EIoG3LDan3I76K/2MDVd7Nk2Uy8mGaExflZ8A9v2I8opo/yIlOC08Jw8P6YKmTid
hrL/J04RQrs/HNFp9oE8nQ8zqObRDk0bzcLha0yO8KRKE9fbUHUXWrK9UEEdBtQq
nwsjPTHgPoxRa/kAeUm9nhAjYl3vzAC7C1aLGfsR9WY1FbLNKybajRcDxTpQ1klE
J5Op5b34+Hr8B8QXDyjHO6Oxdld2+Be8jVb3KDCfcsqM5Gq0d/dUlM2K5aOIoOva
QLS5Y+HKMRAAoP3w4FioUwX79ynetyx1uw2GUfvtHTKG93xhCQK+BD/CXZurVYfy
bJryMRrLa3mOrHw74dj9TRo/La1wHoI8DFZOMn/z/lLjtg9yYtM3zxexQXOFUQXR
bItm24HdLJOo+gr3dqh6hIgOjbAQ8lYWDD4SzKAIur/f0C1saFvUkAs94p4L3cqg
pODdOQFTveKg5/yb3jg8sUA+SAnZWStx4P2gArBWjmtiO7X5rmiBRAJ+CIru3p/A
deFSREmFZ7zBs2ZXkw4QdH/Nn0rfzQdL7ONN5kAaRFt4IzzX6qiVm1ER+FvYb2eM
GA5MMYJdBMKEPPDuJZPaeUCn2Nr9gIkZoCS7DnwYAoExZuHODNrWI/3IyjDfZfXR
hZUuSaqItpWz7XQVX44ZVncZECc5XfBSoAAocw8vlbM1pZxwdS9m3r3dskvHfmih
lZMnhgnW0c7w43aKiS16UvgbHLY2B1OD4hnp6Y3MOcJIIYi9ERhUn1nwjWUMYZjT
aEBZg/D7ThDHWt394gakkWKiKmiqWaMPAhBBqIkeDVyxXAPS2y44hPgIBgTjP0sn
KtY0RcSq2pZCeKehCnv625fxtyBPzbF8gxn7p4oaBKbad71Fw7MpE54zb/pbJd9X
HGgfghCIhN68QOk+hLxlKZHcczyj5bU4V1K+5URl/xYOzxd4/AermjvJMTs2CmHu
3AMLtdXkxFPVZnh3dv7rLYiN2BHZdzX/1A3/qZ23nQ9ZBIT0orKwQmq/I9k+6mBa
sQjnG0KOY4QqehwtOb8w8oP6LDrCE6kjZCFVNb0uGmc486ypwCxnHmTB/bKxxWtw
Lk9EL388h+wA9IM7uB+xxnz4aTMNIZJPgHZ587+8c/o0ru9aa821FZfpCqIo4OsU
j28HWEZBr37j/KgQjQWgOwvDdSNkicOcM7mc/xUbCFd3jzakHAOgzbBEn6EPbbH8
sdBLp/WZTMtv4MZJpaIFYIiSLkLxDliZbTJNveuKcxiMitIdPYyNRTel4lkgP48S
XY4rk7729+HMENLl07rtW95lrjloAHHA4CcWOIYtHDJ7V6gV80rpm5mfVWGtSYaq
NEoFAsxsB3A6bVlQh1Us7OIA9eZuO5QGDpSmBlp9IGPK05mJxrjke8S6Gh6oTtrs
Y/YMkf+uPkQqOTLxU8iiX7euVSiirft0eVQs2u1mpxgmApY96IjeZgMWOTppT3GH
/bpn9Nd7Ke9bHk6hygH98rcgNm0/X5CbjO/wNW3feZ8hMO93O4gKx0EciWzyVfh+
5qFRD9SbJaw5UANacQdXnv5aKu3HZYGfTmH5xc/dIU/DsFF3/KBpzPV5iki9Lsr0
to6O71nKhfHP70POGP+/GBajiEle8GWcV+j/av5CQYsMykR0kTTJLitTsbUqkRLu
fsK9ghOJS2eQCKH/dw0JegHxJlELIMhslZY88Ntr8GOFcRMr2paM0Xmra/K47G5C
VCllOp0i2a4fm2aJdYwERDX+RrIscSK29g0h4fami/+0PCsiQNCNnBzZXRztDPx+
b/nUE3Xjh1diqi4xp2GYWGxkASpH66z+ghxGp/sFxziUfXz2/+8SQJ6OAV/EfMF2
/XG7q3A2BKmehCUuIyo9Dw4LnayOkPFlg/jVoNspM/SFYf+iKEJhbMtoB0NCkceQ
bnvegnIDHMgitC61HVKGNDPI4XvAc9iQAOLXgn1ZK4ptnc/ufUBmKUqag9DVedW9
DVWKBcScgDMUHh/hhzmzdcCfdpQvFmYWNd6YN8Iw/HeBnUa/tp8qulf9PqWzTipl
ZO9XTyxPgTBgJXRlCL1OWCYssd3Sp/65nnYkQjYoV+9zmqV79tOCtcV2vf8q3ftq
frg7xx77ESALAMtsS5vTgzeaHYkwHBX0MeSH+Ea4XQ+oT8EBNI/r1MhvM6WOd0m2
pcgIQeoUQ59vLGGFiUOr4ASKHNWXpS0tJ1WyqLFEHTdjcxVtnkZSPi0XNJS7hz1d
PNvf4YarlvKLOexPyUVVWarkuLwd80iUPpPHI/sUJBG4cLF8swjgDSYLYzzp/v5Z
SgVqvVHLbfNETMfUbdBodv0ybhwtwtbZUML+d6lmmx+yDLryd4APocpKmTi46hpD
F6yfOOK9txfGFIdaxiuUo3vF1YtLmEJA8nS5QYr5lGISw6ES687z53XCqDb2E4bH
ZwjtUuJmBhX6a014CA2WlPeV6cet5cW10L3yqsnIZJ1s3RHnLuRytmyAC5sM4PZn
fRpL5BFBAahiMCZNvhggujyTVv+WS4WpLU6RmVhlufGM175/XPOxIK7KU+CG1Ovn
EXiH8HmNmk56Au7tvrCnnp1MQxpYT77SgbgUTTGMO+x+pMDwyAsImIXxbikSj+sp
eQJEKjJm5ntFV6nSu/fpcDvr5PVQPE79cIyFATsytKgMU9tTckpGsQqQFKUuDFgc
hx3s/ZANH0VQBHKai5tuN7R7oXSCSoFf6wC2f5zP1LTlgLCf7CvlWCODkQrv+R6K
rwwb27YR9xKMMyNm5CviGwJI2YApI/nSx1ExjA0kXCYH+pOn76+Rgow1/PIXy7R5
njFHaigTK8MU2VfgudR/4rd2IyR0Cy6s5UHw6PyyBhsKuppZY4LGZ3j7hfBb4E1m
e1HksPz0Pj8KtX4MkkjcZxAGebuzALYqXTZhqFy9o7keMEqyTHltz3Tt8ivekz7i
uUdASjCtRk+PaK5MJVkNMi+5K+QMt3UNKUuJ8WTmZI5x3vVGDWTccKyxvq1x0WBF
8/TyDtbhZo9TGi5K8BoW5Wjr3p2gHIz75KwQah5BkKfSQG8LcaQD6zfuJFObbvxr
Zvsll9gZzms5OPbL1XyVejp+6/PyYFK4E2rTqNvf8m8MzikG7mS4cOsMZmJFS7bK
pcV27mzlgdhQGJM4r+3AaMP/28QFE05GjisawIcBJ9szi/fjg82NYN5uTZoOLLMI
sfbX0JyRN6kQOoDiKt+RVSjDbCGzxS2o0n3M63NYCa1XjOJXzcTLcwOdZOHf0LMI
bX5qHFAxGsQPvBbDwXE5W/A50nn34Z6Y45+N3qxkr0OqKOO33IGO33x1s88jQtR3
`pragma protect end_protected
