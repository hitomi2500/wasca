// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UJXLgAYYMbB5xpmNlJaG4f2ReHrNA7cdv6wxjYXB4fg8gaTTg0eGUv2yMgejkTIZ60qupJ2ZYaoR
kM281LXBtCHN66qFPwriD4gph9b8pd0/4ZS/fZ6bGqQyE2ojDNchQK/vwyfvGp7/HcezLWOIO6UO
2387pd9ddxT25QyR+d4zT608/ofhmj/NAMf8kxYrZ2KPJlJ7haH5MF/4T4D0SwUMY3B55KPuGAbH
l8jOD8MzzzyVKuiPmgzk33xbOX8Deo9TRPpn3reQMMCeNRLoyzCsMwSUieccBkgLw8O4L8Xe2D9y
tn1KpHc+JjXaheQhKd0LGMYo64HQs4NGZ8o7ZA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
a0Mt9ZtYWOerW5pzY10EnVZyFiKlvApJjUIMdvof0o2Yqp2vi6Nxo4wf+nGTljFp8lGF9gHFy29E
vSwzK+lRVbpKSw1F7FYzFxCMk8mJzPb0b2zz41agrfiPPR1hSi995A3Knd0BzhflwXeNvU3AaK3F
MxKbPlqQd+Vu4bMyKLQPGKI4QjRCUJQ+TTRdASDcuZ20TDyd/WBrM4lcJw8XTsj3pJlboBjeIZ0+
rGXKqfOPu93zkQrZdXw1KKRHPli4ZhQfeI406JemHmUldqjz3dBWcOi04YquFYKCZNh35tBWXbDq
A6+TwSx0arAiKHcekljKNFFk+2NGj5YTFHHpo7fHeGiYvtp8gRnyphIlVygEgfL0t1/wjB8xuIWn
hhO3HoYL0oU3U/SAyyCSbfwLWWlXLKrVGWE3rykOTLB+exYuxmKuYnJSdMXOBHbm/YmGS8ykE2n8
sQ1F2pxvakkzCQlL5qpeOrkxvwGjbbou1Klde5hHjhBBIBQuK2uSZJRbQgshGRnm5pGG547qNKW+
ifjFFLDl0saJiFjxuRMZ8YGHvR8KydwpolQkf+zJ97RvGHAfaePShxBNhx0dnvigReXVfH40MGsN
QjhkE0PJ+MObmCgjrvDc6+NZe++q7qglgClu1YY7PEMWLSI7wfeBoWwPaVvAKoHLqueoZakatxlj
gd2ghAUubEjP0lyk1CAOpTSCro9Z9So+OhzUvlDTuH68ty3kGacaMrdz0mHLiDHMoPhIlu2fgbi8
6EAcdiPfaZVgBVE5MrGaVzvE25nQ7BkscQQcn7Op6KU119sjPgou5PLCf4ClHJ57HAOnk3pukTmD
PtbKH6x3IbNh2j+f7gMYPg9zzKutU+cK5oyfwkLzpyayocEAtN3SlznPhoaLiIA7S1qc8uutdobI
4wV0upQM4FHLRlQcfAZj4+zbHSPVXnqEPg9Cmqjpd7rT9nbIrF06Ur52tUE2rcASgYtOsny7rai4
qTJJi2WA6OAfbLNbC+pvq72af5uo4QQ/OcievSCMENz1svrfbRJo+rLVRFJyDc7LugMk/+uxw3P/
cALUfU42cr5nC6SaMPT1ty/tPJzM4x3z44HJ3me7jege4f2VMO+bKKwPMVH0XZCKYNfAYB4fihF3
oVnrY43bAF6iCo52H4nxMG6dN/8LFLAgPxJrWhI5KsmgvkwWIK0k7NKRy09YlLR5wPOX3kFU4IYZ
HGBhnKXOtvTVFUiJTsIKvLBJVPmRhxsjqnEXgdDbk+KNjUBbydbOVpKKpN1jv3fqZgZzrgFg1vJ4
2qdrDwURIHWKF5yexIc3BiM5QuY7iWmUGUdR/QqkU1olC4/ML8NeTat3ffWIFHfXlGxqKRztSviY
MGRUqubRMWM9sYrd983Bl3SbGdXGOdMzphDfVULBXt0rIZlmgTT2TBv2v8Umyx1RG/X0+zlwBIIt
GCRcNnvs7PWHfVKrkDMK5roiqOK3g+6YZuYd22EnRE9uohHK0AyRbJSOH5oRKiEKgSKIkk+iNATN
e6tTA22x8oDBsvQuVmQiruH3SMXV6VRi2yFtwLwBXpQQlC3+VywEPAfLF9NyQitvZ2Q+K4ffEZQy
vLVGfUhLJojUk9oHgSLXcRH8C8rT+o+g0KS2P02D0Qr10Jv5OPMfe3NPEKwqM/9mi3kphZMmqZq5
WEsK5NyNiUar8MFKe3Mq42QKFWaqTxClvOs6ktXN9TlNAB5S9Z95bWRs0HKc2bi7vwAMZWU8dkBN
v1cP/5Nq5d4lVJ0OXWJlVWLABb7+SaarrYlQXy0YcW1hqOv7GNuVPn9xNVCU2ts8FFFkb6AvjSZB
F4XhkaTaNsPSCVqLykrp86tGO8ez6h4zVw0jGfo/2X9vcbjIB7s9XGr4+6xaZ2o+EcbqvDRj17JZ
PRydPmRDqbLzCmBIV2Hil3C+3UItDG2Jwa0FZEjdkSoGnO6yFU+6HkftLp+o/aLFHK83RablwDav
tb4rtXhLdkcm18actJN/FKHYz7PABIRelXIPnpRYJtSyLiIH8qfhXvMwZW6n6J/Pe+jUJaZcrqRg
KVHSa9ZJcflrX1ZrEa4nI7FUbiBQMNMH7ay+nsK7cNCT7eaDsR9mqfhImF6F+eB99zamUJKYjV16
O58Q7fTlccl+dqvlPViadJyh+IC8aSdfqJs2YfjVpng5+Xee6UenALRieWjD69rWnKxn+EdgP9au
6G16S8m20LslqKCt+3d/6fT8/ZsZ94z+wqI1SM6g0HOZnCgLowsPPuMhGMuMrdZmtrqpVK3j4X12
MnWEhYiMiYPqOSEH0mkky98gTI0+BiD48WqapHprN8F1FazoO7bjfXRMqWcZG9gKWm4POWk2x1je
cbtaEOOg/Z9H45g7BVt+LR7Z8q31aabiyG75pIwWzF5dzznGKyGiPC0iy+T9CvyTpk4VUXGjODoa
2DzPJL4ZWJhY5yu+RpnUGsGZoX41MfNQIpnSHNqcQztoZW07qSEG0E8lPlqIu9fpfgiet/EQ6bIB
YO+tXclHoDSX4HnMuKVCmrIhXgyW6mc35/6z+f+5MG6j4bnu/TpiSlJHC49mx2bqhGTGe4cwz/Fk
J7+IqqCcvk0NZPgSiJxGK9WsQeJi37atfbcq8j4w96r2cH0IZTwy9UekYgIwhYjEnrTEoQ8IBERP
iUcQ1DZ/Xqh17CeNUyXq0wKLzPv8UqQYtaldYWnc2INDlH7/mmlY5IBxyKS4b+v5fT3FM+Ui2dCN
yeDgirc1xh8+wtI7v//80ComSUixCxIiETkIt9EnRyNPKD12HzBnPwlPnRjh/xc2q+zMlRn+USbW
gz42PE0PRNfa3FwUmYc0QqZ+WbBbIaN7BUu2827mrGjocSpAV/G7M5iiqmEtLBiNMLG4darGtVOh
kYenDzUsihdq2lu5NraxyqY+l4oW1L89DWKo3M6XFbsA0jYvsz5BE7yco1ATNUWmtSvBcBaeryfP
GNJgr2CafuktLoDRkIdXmpUaXX4FagKfjzPQU2OI338oB1ZowoQ/0t/PGNUekXExjMXrQIL8BaQu
CY6F8/3shhIRod5NkjWxZm01PiCVBrupzbnjyKQC2seqcMAu51TDK5dYP5fUb9RZtXSJeZHeITkf
N+WxKAdv1AvGt8uhXvE7nUHtB4VrJUc9t9BU6ZPY5dn/jKA/JirlwhNkL224JIFMeq97uIu17tEa
PlaOGck7zmoM7uBFeoXaimXjMq0+67mG9WlMMcOstCDHDshUyO75NnG2B3qIm7lHReCC+fkrEchS
GTLjBwmbUIHHlPjNEwcOelJW2Y6qVJXjRQxyyVDKJVAXk+RgSyjAArHipT1HK6FLXyzthYxUcQnK
hWYsoqy59lYNYHT+bY8yt2t3FE7Dn3P3bsn0BzVS6Q83odi1T5ZUVgVEwRMxUHxDrTPvvgU1lPU1
A96A+GET70CR+Nqq98WJIWbjBSxRM6oel2WPd6MdIkPZYVpr8f7IU7zTqRRmcV0OqLMLxsSlT+K8
xYide7V3Ak2fKW+L8DIjixTwwvnbwdO7KJQW/1EKBaURT3heM+wQ7zrNaH4U8zMIB2ntoI8pw65Z
i8aNnFwoSflFOlrBjcTH/3rjXSldHRDlstILU+bo69nD5OD0605dDVSSrvExXIn3qcGsA/teJqhx
baEFga6tlTq02jNc7iOcLdDqYbORKuk3jHYhJ6oIXcXM4F4oT7jGcMLfhncKH9FHKX/3GIz3/mmM
i2vcPMxVctKfDlttmjrSZSeEz8+nkQAJOlAvac6WfiJjuCkqwie6UhMM3McdwKnJSCzIswQAmjqY
QI5ZBk+iVLJu1c1INtIwZs7Usckc9SqV8ZiTCXHLpIHpSWVdT7uKcVdtaDedVzCFo6GZGyrdJ7Zq
qYliNU1OAVKOlKVRZqt0ZHILFoJVX0jnIs4ifoqFdMbAk7EkoiPZvVlUIGD647LAUptNPcNZBY+p
PwbIMczBo6vqloGXc+Ts6XSgS+iXBsyjUwceiYgd982VgvAGA61JOtbCdrFFAN6TnkvTLYRp0EMy
GiRj279xttMu+u39IhdWRF2rBL3I6EAJs3ZR54bywxN6EySnQ29dA1nXpFWMycmpWSjZOIflTUkh
pjFytRGxI1rGUt3UE5px4IX93lfmGri4QTv1HpZPtql9r3Qgb/MNlwfjPuqAk8JlQDycIl1bkevQ
3Q80Q+aPYJSoS0+TGba6z7VXZNdsCOj1ThLoAaVX2nGWk+ZvPhz6frBMPB5snFJTC1LdfF+gwUI1
16S0a0Cnlp7vwN8UJsVLnLXBjCHgzpcTZ4Hmr6y2plvy0pov/VRumG5yVUqRkS4pVd08udJyAzO+
f6ILHBnCdEJND4Rl2C3CoFWW1ZgnIMhlMzBAajQq5Dr/xBeOTdySG2+kjYLkhJZxiNJGljDP+sP4
q433sERXtwZQ7IrZD9hrV/rlwGtFECDjXVnFGVxV810dwuyl/U0lZMiTva0utGLGNQsSZ9PwwQRO
Qcs+qM58FLY0wDHWErsvNvB5fgO8uUDdW3ze5Xs0n6M58+oiSpfk3DTjmIHizVZIUT2g4EMnusgL
7SbPokP6w+1YIAF0roUhvU8XXLk+/Npw8aqkk4myYHSaFp4vnBHi1C39ybKajDXggBYqDT8zINPb
eOZW4gjZW22+V/I8x8EPhvu/vAcGj2Mnql3N+dnEvr9jHGZgjy5QNGw64KLhyKCRkJoylT/3Z83T
0PqSx30E0ejJ8kKNogY8k/B9syRdwyDPKniMK0k2GEdPwGesvydg8L+mZf1M2t1aOwiS/YqONX1L
7qUBYbCvLUbfppqP1kDtIJ7httBSlUmQUxbC5Y7brP6pC25alGgG3ZQoQmCfQaKUtFz8saYuJLU8
QUezC67hlQR1SwDIDxGSx12bNy4SwfjLUj8GMjLCJNgaMO/1oyjjtFIQXGoNwbJ0qdOoU7TcygZU
921bbK5cbAMwu+U8BTXPRpO6J4Awt6rXSHa5tyjtp2GaoEOwjqffhgaBrXZaWZW5btCnzTkL7Q98
Le+gGnGLlMd6j/jlFZdWhPhSpTgIKhyyWdOGSZoOthzlGeknXXZdqen/wuFa146qet5LWBxbcr8E
LS/EQj4YsqG6xCFj+HFMCso/btr+uBiCBqVZBn8MSMhJyCss5ygXAGJ0P8qmROBfMOW6lTx6K0Jf
k3xrM4RD0VnNncFeQPumlWB6ABQEotp58zUVrBgu1pBzODQ8vbrBDkLJO0YHFrIWEx5wP7kkcpjf
eNApIkWXC+MRniGgJZqwGukxRSyGEAXw1Zcs01x8x913+RZvz9ilQCJXnasDlLgNlKLTmyJ1/QCO
NzyrjAeZYWm8C8BIt8LQIvYLH98nVomCWUfJMlZ6cE+mUIxfqZRVxe0rldas7KoVX4mfkk1FS0o+
IuV2+mv0mZgj4fuaHdoLePTXjJJ+UkabWqppYgwIjFC719KaUd6neYsrygomC9aEqu7xuPmU9w91
VDXV7kBIkBYPG3b+krufRnRkn29oqkjSRVsupKEHXpyu/V+P6XxgUBu6G2ek3VDroWLdJtXGG1Rr
svalJAdIiADMSphg6We9VyjhxhTCA/qGUuLDyrPfSHJGEciB46Wilxz+bIEJSXj0TqqKZRo3RNWl
+4m+RFN4RT92BRYHTGjtGkyr2GU30HYM0GAu0uK0gIQNkb6ChYhJnPWOTWIlssOwtwBil0rPng9V
ZliMpIwBFXHODpn9dU2lEmy9iVkgkAqTWws2oX+2NGK99+5Saz0FMdJkp8B9m9RaycYUBPocbdvA
ZN8+8cvkI+r/t1xhOVhZkxHHUW8HTXp3NspkgZhfeeh3XwEVJDubYYc5MVWaVNeZDJKlQayT1V8i
HT8PbkzogZCyWPQVM45CDckyyLNNW4zkiEt4Qeu/yRAuZVm5SEWHLSbAMzRK1ARgIJ8q2n65pgbu
e7q82LqdRl52WUvLRtwm5EZOMLvhmSJ3SzfEkmzO0s2bPPleYvqi/21QwcJHVdhNTjcERi5mXHMh
RW10COFKth5qTut9ppcw7lcpxdNBHINkP7NbP7y1yVvZwm17P9AW3tPYGKnufxsoibbgKahPEqgl
KShpeccYLR3PBP0tOl32ZyltyL+krc3xaEAQT8a5O+zB33ptMlyLEX7kcftlhz09gRuX9UHh3wcN
G4QE3QVz88t0DULX4Pw8MN1/A9Rrm9ZTelMwnZVHrEt9PJn9lrXng83dZ42IUeyJ/IViEqwm3Ulm
0QI7umS27o01PYwh9xahTENLIE4zIE0FKJ86fY1YsnZnzk1MIe8DEDOaatF7y+f7M8PkJgUyhPwc
teyioJyjBrQ2ONSU5HAUR9rdEKjpJeiXns6MPUX9SNhL6ub2wG7N4GFsqdAaHcnaThfXa8FCMWOT
AaACjtdbt9gGPyywzM8gA1miScoBrr9OmGGzZol+nB0HyjKyLUKmp3tTfe9nWWaLalRI0Y5V5nEN
oTEO/stkIivJ86YU2r0VFQ4u+tjQ+3AiK6UTRFP0PF515b7BMy6D6iyn62iFACWw4jSb7w/e6+Qi
B8rI3crMSPmpF4TxY0whTKxs2SgLPU2WPxxjZs4vZbIDmXtLBQok1SoSumcd4e76r5ApQJzcHU5x
ImXFLfSwgkjhxt3UiUr3uTUJllWnAYQtD1lSorMZ0teXTj/m9PWm2n32yCB5Ks9vGcIMJGeqtJO7
kD4OTk1vjgYl2I2JPjPiWtP9+/3m6NETgRcTVnJWuxtK6zrY29hI7PcCatKshyb1eJwjHJi3EeYm
2o5oRjvMSipdRsuvtDGkXMcyVAjFPHSCaR8KTTk9OljxJkfg3O0qHYnRHy62MvBdOtxPCdYMQDgQ
CZ62Q2neTgBbl7jAhxe2pKtXbT7nJNDVl8DN86JHSp0ZGoS1uY/5h8JEWGUR5iRruBNUdQME+ZXq
T7ZZHivh5knyWdFdT6g/rHkhhjyVSiE11a/vWwwMXwvPmltEHkjKAgmCTdKS+o5eQKKv3+SO7FTX
ILpMcBwy5NN1xRKCfJeTTvDqP6CDPR+WiJxijvjE/7NXNZja8v5l2lCTurUiMDVadSU22jfwpoNS
nRD7jjKwy5bpu401AexWQub8GVUGW3scGoZ7ZJd+mjL8H80y9mcmED1bSJqIwPsB3TTiyqwrdOLp
/XmsHt/Y3ffhoND54HF1/IxSiiyt1WX7MGRw+fDbN1rpTVv4wW3E8G0FpcspWGKRy9UcJU2uL2tv
q59lGmnRLh2T4ljEmRCy+HNNfpydwseL8xpx4oQ4azBDGwVdFcHhusAkTbmbGJlunSyg35E8ID+h
1eYs1AQtl++8o1xS4DwZhpeQoQ9/KA/jE48VO1MNBMgqQw5j1pkf00WQkj4hSdi1Gs8S0R5vOvqX
kSygFUCwXhUv5FxKQD0Ljr8ujbKEpnR8hD0DnCJusO1GtN2r42xD3OtQ7vzIyRGYlJgfaR3MnT2J
jdOOa9e9O1xlmN3nTkEUDUhbm9T+eh/csol3+/61ztYtKULJSXlXnMC3T7i4F51LLpB/y3Iga99B
XxaKUpjiAq62bRPrkjmFaBmdAU27Y+TVUsrKD8YGyu5yvJFfwbc1s0eXC933E0MTDC7CmD5oTESU
p9LqIOmKkhKwQgSf9PeTmfKc74yru8dp0od44ZtlRdai9aez1aY0jTBtubYweQZuT8J0W6BZXe82
st+WSzUb9rFQz22ATXGMaddx8KDGNM3oBJVD84aj9Ucv0pwY2zHGVuHTDcciSF4GjWxiGBuI4bsT
c+YmG0APRyhKK9YeCkdfKxBXoW2HKpbH96+Ebs30LR/98nw1ZqavOSq6iH+OTN3IdtktBGKB/ynn
7q27zPsdboaEGKrnpppdVpjeQm1UP1aIebQ8viepTJwgVpm0krvLll6e5RKSbYil6c18MX0jPImC
6uLWq3NC3Vekwa6G3T2aOyywgURmFX9Rjs+tJ7L+dTUBGM3nnS+3knQ2j1BtEHx645PZyMv7007K
Cj0RTURU3iwZ5nW7Tg9sueeOBJ6ixdQT3dzXnkuCFRbVXZ1Ha7ywxShBHSbairzrgUi3Gp6GGrbT
NC2vpckajQaBMU6OrMqEsifukTflHlFnHJg2UbYpn5EC7h16Sec+RDA4fnQiuB6OJsAz3HskzkyR
3kmVQmt7gI/pQxINwJ7/rtXqXITVnzzKXzKtUt3aqtGq8JVkwz7B+B7qgDaGA2ODs7t7gVyOzcIv
pNOnlsisg4Kzu0f0GLvamEOCJiuQzgMmpwUXkSNUJW5kLqCaeF50tNVNt9IKiOsAtiMWUkHE5r1a
HjvyoDTTCYLGEBiup8I7YtFS5keB/oWzDvoRpdK3YJpfGqBAPd3QEF3vpSEiPXqfInLEWpfObK/D
LQL5lTsw6f3/DxnynRlD+KZnBvqWJhN2byDZDCpqT++eiQP7YDE/4svSdgONjv/isqqGBEtj/pCj
V8qrVXu+jYlOT0BYUDmkxUcOTpu+Djf0rF9ypTiHZjft463JJqfCtlHV9vT9YPOYRHglXpu2Sup0
MFS29IASBGuUdYnIeibDmQ29jzQ1b50QMyBVKdtxlZ5nkQ/MOgb/CD8gNR1YcHlJ1F1wTSaTwwT3
ey60XUt1v1qTGWcztGv+iCwjwBY+zHmJw55W8apqVrPMY1JotTXvV40btVD2tkooQPCeu9x5qnT1
dV/ACK8+S+6E4Z42G1MOkSkpW7FIHc5GOvgs987O+3E5GvnyWbZ1vKoFnA8Fe2JjcmdamvLjPUG2
PMHPKeBqCGjTe1UW096JM4JLgzcDJJk1ioNaVyffe9WVt1+slnvI/CGQ4Tvn8cllTsP+/A9hK3qS
PoQoafX5WbVI4TSd1/izqW7J0Oq6qGKXJostwbCX2/A4hgm3g4ZQGpu24Dc1Ii4Etuh/kLW3XNWI
5t2a4+Yikg50f8EV/QUekOK8uueXmndb70b1IDf3HEVFxdZI0Pfiso100X38tOXSW1KW4X8HxFuW
BnrISgqPy3MOSAy2U3VviM6F3LpGhVcdJY7hXjn9gG3meei/hXMKhCr+M60XMsJI/QVCsZ8d7D+a
4z8QrUXgFlJkaw3P4MIR9EHEHqseFFDTIlt+MzX9LmdRBjEtxcqqkDjviq/K1Hooqgj19e9y9U8l
NDB5TcOr2UzTJ665td3QscdMqGsln6JbAfM6e/u3Td/9BDGLQpqT8PtPYshGGtoC1CXSbvMQsKul
eALiiqd/5r4NcItfmRuNY41maXVsjlHWaFVpBoscb4OizJc8TmD2z8Suad4z03wxoMQU+bMfgn+s
HxxpRA0eRh4MiP1TZnTALIrCmo7hL43YCrWhbvPGrV1UjOKfep71dMJ5GhDkC+fvzflm81xm0RD7
RYcjer/xCL0ht/wcmwaLcdMaF/FxTCzeA8sXbIqRXHyvFDv3y9KhDZIGbwMP5mnVR+T3Ah80cf4H
NqqtLI0Y0ShfZpXOSxK5ZhUOIR4mPY1kkmyt0+IfDohB/GI2QMtYOUynHLSXpAsxs5sm+9TAdVv4
2YMzvXYkC7Mi+cxX408cU1j2nUKa3wN+jW+YW7uTV0PaNeh/CgX+MpLgIXTe/IhXME/H+l/IKSSo
SdFhnSAn6Ld9q/324SjQ6DoLkhGbLJvHR8P/kTytvX9KpduJLGJGvIoDDC65dCUvS9MAHjV382Db
ZWmiazavikKtyOcTsJpVkQGJtXRxNTahmsAJAhzLC7Dkj5OQFdvqpLe066TM8z8IR9Gdgg3yuLxF
v+BA6wtvpNPL3sduAYLghVT+dT6T0oC2jk9SIOnoS49XnZ7iUNxWdN6UDP21rNyFzE1/pf0d0l4p
JccnQyOGoutm00viRH2pKDsmQaE1bFSPH3y+nU/qucr0WEveLTtGmYYjtToU9SEyHJqcKo9rYH43
dGNRh/EHcJBtFOuO/+Xrk3qC0PKUTrof105OqetCx3a59E68gOlNfRN7OZURypnWkD9+MjzdCWpj
E+/cI5AJOqbnn2YJmdVtPqSXL5+Q30KFrjIrMSOwG/VPwNswuBWP4hWFuhXboXI7gf7tH9msH7Ki
khPq4/lTjCJRLW4XYSi1v5lpM6/aBKco+gPXaKY5s1mrSYAEQk0WF91a62p7eLTG7RLgaeCEptU0
XUC0R/h/KOJq8aezwoUyLO/8RDoT7ktMmUMu09eP8/1O4Vv9GnexMVH6SH8r/w0ud8X59g2FGGBL
COjtWS6hvmKuZNCcayoYreF+jT7EqLVTSPyuXHg5cJXgMep8x+yoS3onvaz6FQHAhSFTwSiVujeU
Bj6vm45s35Z6S2ldWrYbNWKDVEbnx+wFeZcCj9biw1tnnlsdvNlnnl8rKKcb9/191gZPGEv3jqLD
5AtSAWbD/FBYiIuo1fo2jY1GX3PnmMSEkROeU4Ju7yqWiHzpNQvWFGDYL0/sIrsCwPy1D+74ZI2J
sX8El6H8Rx8Y4z9gkp+nZDhAeYxBlatFHGJws99ty1b7awFczTMe8DlACNrKzi7xMHgzcNzW8aAM
mCesf2v/QFYfgncMln9D0oJA82q3ohW5IoWpM8DjXoHQ4QqYmvutrB5foIIGHcuxjHgUvwA8NHHi
Fj9+D2275dp3h6EdXMB7dyuaYlIeE5o3HiSKr3WGcGNyhYK3NtM767Uenjc3xpfsl2s8MNnEM8rX
QS0WhnGFCAWG/zYl/MhUjWurmR2akOLQ4QASWiQ3tde9kEYn0pOE2Yn1+1L7NnFpZGMsAOZcH27N
/wYzFIVdiygWIy+CkJ4v0oM2RQTIeh83OxE5zY+bQVN6Ra3j+DxqwzuadypRf2UvFZlWKmlgtz/v
RcXWtn3IN4VV62YIetI7qCQ4fwm/b1FATioR0Os+lmReHGx3xMUmtx4e0bIGRVA0sZxwnxJcjsjN
/JnwnA+fb9Uvyxlsw5bgZ06cD7aN3tz1gg+uOD3ATc4AAQsYTjKGdWhMQiNepWdp86nq4nGnizGn
hqBI0g1kOnfHtRQ2TPsLmYW/rwxM1R77lMS1Kxmz1WLs4A1CAO2kFLnJtJ7UMHUwPMvKNoaGiRhL
y4Gdy98kGy5WxjtMrfoUV8FFl1OnKDIEMWjtuk0hQEWYcn2mIPhMi9SFcW3LsEq524MmF7FQHAAx
1BjHmQx3n3VtjqrgGYXRUU8LslR3OQMW2ojpEBZLmTsEujsP7l3mLK1JC5UaVt/5xuhiMm7ViX73
fNbNn7YojTBW0k43Q9P9E64zRGCUPXT8GbTVhhf+h8oyyZqaStuiZPgPDnSMKbRdx9HGZokOJ5pG
U5jUWhDVtMycMi4AgFxddMruR74EAQiiugYJSPot+C1tGrBoSDDoZKDsd8JlduaUdDdi2i9zkPeJ
KT2yHgnuOQQM8Ss14Puigp0D3K5zFReFGx6q/mUw1gh/BDkALCEfGoF/i5qz6cdLz7eDggQhMsJ1
/DMH1US1CrNA5AMKPN5mE4jiTlX2U/4Hx2g7hkXkEtvOVVbr8IcDvJjC2Ds+djfjv5ewK8elqj5j
687aY9xTYeqxe8Pzwr6pdtLp5UXPLOjxCN1Hn7/F39hUVlJKVFsVu0iAcJCpV8JmKB6ltzgrLOkQ
1TRSbosDt6I5+j4EZLASK7MuUL1Pkjg2Y6/jLzk9XaUIo0LuiEyaRBRo6mjild+2TgbBESXtHgi1
LCzECzPI1sSfKIzUB30EuHtyJCQEQC6j8/Ga9XmWHtY541hWdgcKfNmJXvKy5j/nszbYhiyLVcol
GgdnuQOUf6x8o+Ej6prBwY4gueKO4eafVhJ/GFT7br/JTpFtWkPeDonV8y8Z6rgZcK/XnR61fHuN
xGRZydfGHzElD9I+xC+S/AolOrjC+VZmLadBqBMAMdmxyz4bmkcgiQH9d+MtXTd3qnm0eXVLA+5u
C128Q6h3ZcZtvJ2SPF3L5xuFTBveU5XP9o3JBZt75ViySpoWlPkYvpM1g1LQCT8uNtLpa3mcAt33
PEo8uwQz6HgUekTmn3sCHE8xaCOsNF/O7biABXhpVEkMOznPKbuXPCi31EWA8fuAZYIyBrugC0Eg
3S1rxVSg82DAZLs9H+4+XWw1KBaBSrUGKVa5sqPjdeQDqnR5rx9K9Ga83NobxehhjBNJty+jsOEI
xkV2FStShUNTrMOetknnKFbjFyNwBX/wNPzx+kgqT9orzxpdpMCX/963oGGPMq8HaCpAQlYzF6lH
/1GPCaCXdRE9FxVF6mgXZfvxAI7znzhILrgKqlkQxGekIDzSqK3z1kHhWNBMJ1hz4wJK8OknEGlk
gtYls1FY2YR6bdxhR0sIDBuw+ZyKZ9PmyNPQyBtwJ0wnC7jxkfgS8oaK7NxvRkrx7UboBDX/1Rsb
KECr2yGz31sRUIicwGT45pNcnLdkl9Fn566oRWT0nH3cdPIQZvgMztbx0b71Qw/JXsDKjfIaFiYO
5uFkMJ/rq0eh9PhEWmYUigdkJVKH0KojXHumbunz35dg2ixRoR5JDxOkdTNffdEG5A9FF3we5+Ix
5aeHC+9eHNjCVeY3hBPnkLvqs/WFfcI/mY1t7W8AV9EoK1yPNiYFbGQhsuI0l7UOGOAsSt3YEeQ/
ApgF6fIq+uMoJX7/zHahFg+89HLLYV5lheiXnnCOPS+4xuCJjynzvEirYjuedZsnaXHQS67extnL
7LoppJRu4vCzgMZVU+Kauis64I+QDVO7KVo3QHRyd2JfrQQcrno036iWUP3vt1qooaa+rwPQ3/VB
sDJw3PHH23HMy48km40hFVuR6fVutA60ErYRTsH12g066GO+ifcRNZipoCcZpFyxvIyg5vpz4w1y
AENr2uhri8ZKFRRrqRuuMFdkDgEj7RfXqb3jDz7DbJ2AeK1PHbYGqLpYVdhc9Km1e503KhUY/tr/
g1IYpWy3u8tPY2HH8T0padt85zFfajW+aDWCEfGcFP7FvjqYAWyWAYWkRdLCXciyWRk6qoLtsNrP
+qCvWE2w9y2pgBYq2shpreBu/Fy8WjLumQNlmplXLt2b61H1NkTk+HD8OjelZ5l7wDgev8eo65eN
s92adtUak6Q2Mzhq7XPS8N+vav4AzHyb34HOLiLzoTtFJaJwvbqg1cuTbuLTUywKCdIXNkpaG+mG
u2GUgW3uIkEtz89Xr5UtgSLiuZXf8HZKi6uqsCAI7MWbyMNWzL8Xkjjy8WjYol8uMXtT7A3jnIaT
3T1nRZt8LBKikV9p+pSdbm3WQlcK45OmAu5CJspPT/vYx90z0rmHgcQT0h7/uM6ypHmlIiH+iJgp
eF9ED6LDbQITQvXbV/q9ooayTXUCDQ2zhrpZhxDRQvEpVYgE+bkgXren5pcayLFMrgst/mmhaDEv
kg/kZiAP1miXS4QooVExOQvEvh84SWxQsi206rM7bk2cr+VIW1Kpa3/TVCwWw9Ru5ttTmj6blUox
hga22mqwsR3d6BO9W+y6rHHmexAVwN94TL9k01zdXIE4V9l4lkFNuALCXMlWSuFHlHxYSxyzVqGg
1NtKPC2IjISA4Dx4ygIKlC7unSTYXEksDjslAIK8zm90KyTw/9z284dhAndRu23f9fRKRN3wDFEt
BMpCOQzE8h8QuFnL1SiJURf46i5YOCy0WhsenqhZosCYj5dKLI3468O+2DG75KGoFnWMeY72QNUZ
vQyyjjUDbT2t43d6ZP+AiBQMlYRs3PnIaLlkurF0axf2KU/2ELk1OPrX18mQCXb6A7BG8ZsLBuZP
WOFMTUrZQxT6Yc4pd1YmsimDsOFt+vkD6M+My0HZyRsx/0IA6T5yCNMY6ld7ZSYULwmP1Dra/Pn5
srBPPi/Wc2QDltBVyuhD+OpFsilO7y2mQxBYceFlOrV8vhZqppcUAM93SsJlyeefoAHyDuM0IrPi
CwYC8gDbCdCdOtYYuBphlZIPb5NvIp4Mc39XxVp6nvIdHSzkLy1OJhSEj9tMl9p2gyPFknL6Vkxt
7j8JPldiRD7k423knss1BZhzojWd8BnXApCOePZPNK0X25dTsXzD/qjHh8O2fEzsarfZamDixC/G
QlR9tZFS9NpRD/aN9QfcGZ1Ps/LUPxd5FMmPr5JqilCjkzQS0ovG9Mp9z1iUn58SJxkPvvl9Q1hI
ns9iS+KsLVXMMWP4LL27PYbmCpMPG/UXU+jLeyJMyko5c8shjx8y2MD8+0vou/I9g+fU8e3INoLl
QmL1Fdv9hqg1wZqyzcaFPhUuK3bTGpNPTt+kLSoKRYctXFFBYTKS3kIyoGSEc2uO3wkZOmlKudcm
/ksMc/kbqG02q+vVahbBKfJCM0f6nUHOstZT+QDX/3pu0DKhUVWbiTMBytZbJtx4I0bM9gBxXFsb
09SKoVqtVA8uDzDmuoG/ZPbp7Qs/536dV5ptU884Psz1HGMreLnq4Fs1eUCojwleWIYoMRoCacip
fFm0L+ya0hG55/H48nAPx0E6U6f1WgCweq+/vEqxXpjXtvK0CdPwxyrfukAt9B9574XvJC+Hp/fK
iEiUKRvi3+sozIVD9oLaOXdpT4QAJecska9EFILB332wAl56jYHzIVoOOt7AZkbPNsbGWYSB5cy3
GmQyBiNJTLr4KV3AstIshHp9XW1Ur2uO0mwJmySmWDu/hEgVnnl1lS/ce+iodXxKTdDPm3oKPTLO
kTCA+rT3S4jonOqgKm5QGuTyvf9MXWluh0DSvuh0tgnWFD6fGcKCbklDS54b6i4QtTM4KAyx+d7F
Ngco60FJg9oUZwB2yM0T7B0O3/9nfz9Z2Xa5eqnT+9zZFX2garA7jFPiOgl13pjFLxuiO+xa+rqs
YglT0tzu+H7wvCuRoFTUwxh7DWuoZ/gHU1qGgSQ/UB5FmQ2vfd1FVSryWFQvkC7f09oOG+LBPkAf
nlKVsZj1zjORHwV7j3mGLaoLA2cetSh8YDbJM0/K8EHCwGJ7sWYUjLk8JZOQwmRFhzqIkTZmdAXW
CPDBmzenu+8z/X9tdRaQC+kbAW9NhBL7IlAjB95i2eU8Y5zwxP5+dYClQ3Em3fO+ou0cT9uwT1uS
5CccipXKo40Z+jjLIzruBFiA6i+qu8Y9FsGvSSmPsfzw9FTxeqkYLz/YPmh25o+VTSe/b3CSnqsM
AVodLqwma383gBAGGKIS2NcfCsgcS9CWI7V7egh+5HqFl5fBPseEJZG2PiL//Oa+yExi2hzzejLQ
NbVeXHECHzydWTOLUaG7eLL1BpZNL6UsXS0QbHAAOjXK6Ab8/IwTdPSVlPJXhz1Ufg2bRzgCBRGS
9HbA4NPirOKxNwisSz6GaMUEM5pmHRYvXzjsE/5ZSYZbdvHl+VqhLhblFpXuFmQM4NaGK+ea1jPj
/dwEwCL83WIEi3vgCDFaGSQGEFvJihhLVjOtQpnEyNKC5FNyBn/A8S2WN4FMYw3Y3SWuOylntSPI
PwgyBYmT+S88RbFit86igHjBYzAkqhhs3GcI9IM/JLBG76G5002koZaomK1rVq8oisX+k8HYVp04
saOVzoYV7MVCAO8XgMtaMrwCyN5yrP6K68A2VtV6pYtJSFTfI974a18GlaAdbjhpH4xLYShLkt7m
0hSKkQ==
`pragma protect end_protected
