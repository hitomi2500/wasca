// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U1g7EI7rn43t0ndqDFTvn+1Mi2/UCYrLSVlNG92Qs3/hI+GwkhSri4hXGM1v1hr/
+Bcftj8TihmZRfrng7OcNYr+DRniaMADIJYVLvLE6U3/zr1GreSUqG0BjgNqi6Eb
EVPsdyKEQwQrK/6cVTY0a2P68Rs5u5zi4TT7vXrlCKY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48960)
YdVlde5DHA8YnBHlMcO7WRXprPA/QAreq9kloVmV5uk1f0WgXrOv+zHKheazy2++
0E4BB/t/q/0vXdzvDDiWoL7uwpoEhElggfIsoChUA756ey4+fAFJLdBueRyNqQ13
JWPF6s3vl9I5zNL6x5SVQD0CqJxdDSrBAv/j4EW6Q8Ho7TsENYoWoSYtlYbTXpNs
xswk5jU1BjVorkDVghTJ2agFt3HPC3eY8v+T8Kwp1hUvp3pycPUjqJIwfuxw694j
mIKXXMWinzmR8OVKoFQRuv9wbY6YdbsuD/0UStxOgzJcJ9HJaJ+QgwH8fdHNqqrf
6g5kN5Nx6vcDm0Zts+9BcPDI0Y6ZGwlQAAxFai73A/j5+K7km+1ZktE4ZGN/+PdU
/XSdR2EOeqQUTyAyIrAzS0oxLvlVmeksv8JcVO7DkOq4Jw/q2EV/JMNKL+8IDJpK
zcW8w4Y2KBftWMAU9CUk4wrD+y/IXEstfG0m9Cgxu8ZXR1ajLwr8XprtPWCqUdCg
FaIjmg+sZaeMdjo8EDtqv2yn44QntujmY8Mcl4tsdesYOuCArPNeGGNfVDG3ikRP
tQxWqKkcoYUNQtbfgkMWfPFUmL+DJ990dprcBJc8YIH6vZuaoV0m9fEys/c8Yhhs
DLzeRxSRGcK0FzjPxi/0ArBvQlpJltUOV8icUlXfGzDRuT9I/3jJBJGKfcTjlBzE
+5nzAYkWnFB9YPsd04B5MacUn04o38hawiW6mHaezhPyrM/wRwVdX07tbspgYhbP
GSFHyIt/PJ+rg72rYAzkF5HMiHKQNeqgagj20PXZS9uBBbIQlgVGVhUIFnghCsN/
5CDR7c6uX4kTFpBniVdxFdsB0Jl8zt+9221kme70jNrMZInPeiGS4IxnMmfnDaR4
3FTNLOf9CNawR/a7ur6DWNDElg8ouE1574QSqDAAOBMyf1hwhbRjQIfBEDTHfGqX
TK4Hd4BpDLgyMPweA8KXs1ubyJhYNk+dPmjhJvQc5B/f4qen8A4sYog1i6tXLsNO
nhMHUDpx/pA6VKRqvqNzbRqNlPQ/lhizMtangiig7RYfiq14gMdXOM+ut07rUj/8
BB40PM2KXsLwFz0b3Y/Vm++bFxghOvJBzCR4UmJDXgOy2vlF471ptY6KNPFryE8r
NlRQDaaSZDG2XJ7AtEEyblYZlQjCWq95fpyRg28VgYU1DyU0CfUO1ses8eH+cbfP
K5TFtnfAXyp8ZF7YA7Ay1Lwnf0Y9Cb4myGK15lgKNVC6/n2SYzYVznVL4gAXcgl0
oXwXio0RvRVnhRFruYEwcTU+ecWS+qptonxDIWc8pQJJAn8ZikmToV+0upd5xmmP
MxdnXH3xq3DAX8TZaKruT/k7CVGYVkEllSsizb+aHQkDAfZgWKEiGVXp3UeRRIoh
aiYCyAQgbo2rqNltCM+o7ltLJY4AQH09a+ATh/upby2WyreK69UJ7DlSdW0IB0hA
2Wul3xTMktIXoHmzJZ8Y+YpzKmdiaWA6j93dJbcU5PxAVFbO5SLdeLzd/gz7HUyz
zZhfDz8E56R3Yfk2sLWEti/g5I2xX+OoXWVv93BZ4x6Lbc3OjNZUQGl75ezLw+sI
AMbUhSrKc9QpUoE1vjnjXo8bzWiRVzPM4QCJvVHS31NUovoKhckORPNOj5F3R2Vy
zEy3Yb767kHWUCrHO8UXNRJPSLfGS1F+r8n4213My4He4VwHFEqbhilJbjmyIag8
usZi3OGXy+4i66bfgWpmSGVQFncV3uYILdbZjqz3h6zmwOlKuaYYrTPZvBaGaD4M
qbqpLN9Z9OnmFIdybY/eIgFYuYUIpSNVJJpWipSi8iI6g2J08h24MkQETRN7RdI3
9mmCY/vm+0pbkaDXtb3f66HfIFeuWk1EzDNmObu9RE8i7U1idHj9f7XSZ89TgaJx
aiCIVMd9kLbKXeCupGjsz5B/F6iYMP2HMkX2gaH78uMxjB2mOpjTi8TzdqiILclz
eahiINevXK3CWrHRE/dfR+OBFiQNYpyFBztnHMzf155JhNcRkXzReVt6eGjdGX9Q
i1tDCUS6khb1AUi8ZVcvXRhTNw0cQ6aBXjAXAAUVuZYbGL+PyUSxfQpdzWnUnWfr
WyxelWMruRR9A3TqJatTWtPyaTxAc2KIWuI2fIpqO3qcLcb03xyP5F3jMp8oeTTp
WXToiFqJpf0mStNi1FurtjkqMSRK5LFLlBgTqklRAqKwslAvbXBUi0IXnz1Bi4g1
PbsMj6/KlY4zaiUISw1njPFGocNWGn99Y2v3VTGrf5UjrnHReQu6LaR5wpoOBfth
JHr+1PL6mMVWG2drYxlS+Cp1MHsVpwE//q5V4K5IFzSnIeT+L6nad6WdtE9igMe9
r0dK+gioV8TrCMBf+0YwI19bwJiQAy3wqrVxIlAGjZK7EeSqSx9bMI3MDWhwTIt8
bGaUYOWHHd/coiAJfatcjHkxeZxfGWiFOCRLWe6zTrO1TobPG9Arw3bZ5GZtltUU
BB8t/iB9zYMatPNFn8/1ZhptIdJ4fpt+xl6I08cNvtzOwJ8EzVn192ubxaypz5nd
czbYAw4b0EECM52BfQf3gW7QAJ3016XlmfwF2iF12QmreD31f4fp4bCPA61kH3W7
a5tP3EEWn5g1iPkh74eO6QQGxnEIHqqugEi/0RKOO+PU7AEAQpGfj2bQAh3G6h48
k07etUHGxn64yFmpMx2t5i5FHDjK/uBaYRT7PVqSQVGHSuB2QYsOyF9O0udo/eGT
JRg7+DYQszm0uYqhd73WUT3SiGKmppnwXsn3bTrdyTn/nN4Y+XkCvwj4BXW40ivl
bMznnz3Hefe1t0Oqk2A3amGiCbUfOa1qJLpKBE6U81OSKwdRrmO/x7hKBhv9hd10
jzwWAFOHqfTn4RILEpFeX4E7w9Z8FxAm5bTOR2fgAU9ASnYFAu9apQV4DtpK4wQS
bLMsLZGNbPpgn/gpTXdCZ+tc2b/E11buyx7CTwSmH2I3OGt14mgFV88Z9VdKkWnY
VylRGkTgkA046kZWTl7CYKjdiU7o71sULpssfzJM50Rh+CJyAFofZEaEafdE4jGT
zySl1vZeMxrC/I7nQF27MAHSndn0NdRY50JhbdpTB75pjE6CYEqmni9ttQxxAZYS
T6dpbBfNxATcZ80F0nYuMgw4O+iJflYMSgZNYM34CQ7SD+5kirnW4bVr8jdlfkVc
uASagF45b4NW1gwyp7BQZz8npLkrAUiszIo5XoOk6/lOr0a1etMqcH3G+DNiC9pg
vc9YerfCY+rDBjSd7bVvCCp5cY/nzmbWC6aZgR8+nsIPZT9wy7OO/FAX1vyZhfW5
BsbQqzGBmdTxkQGduTyIalvQDf7jjXboYRd8G0/eMltJH8hSoCiTZX908r3v22pP
n/q813B16cbYsfxnd/5ZwgeTemVNQO0Q6dsX1IDqMAfbcdM7ZcCUYKoD88EtqpNp
KOSxlTBpU5clT61Arn/jnTuxZGR5V4c2Tnq7KWjkzbPTkJ1V3CKEX/CCXHI9HnJk
PmFjDhUXEoBrdB5s1hWpo7yXyHMtJoVAu1+sbNvfFtvmBxRfCSm7NcJig3L7YJf/
Db2UFcn38sdVUZYqGyGEFOrDaiQ0cXk4gTjKLjc/gdb4ZAC2+gqtry4L39sTC7zx
0MLmC9gxIydRfcQLHBJDrnedwzGajOAhO8+Y0qAyLTtLN+Ps7E6e82ECG6xepMUT
bQIM67COxW07H9wakKti2UFeyRSnF58DLclMqtWGm6deiFZstVA5AE4uCfXlBPBL
8ve6hZfoY6RGFHJo07gC8dKVpWt8HRs29nHbzcdwg6deDgFe1XBWEd9we2up1XHP
bALrwBpCDKzEouHCGMlhEYacIzu22X5WPbqrQt7p3thEYyKdD4ePGJjpW4dIntQG
l7tz0ibKcwGa9XwPx33SSqO4a7XAMqZT7yegmYFfAiGeacbr32cZrKQz84rKSN65
qmdTa078LBmOiEdSSt2QYCW8AKzu63nCPvQFltgNncPWTcR3GIU4MklECZ+LWl9A
NkA4+Qd3RfCogKZyEGJ4UjKbiS5BykalS+DeLuu4nAkRwGXCRhB6hd0YWnw8w3Zs
G/EUjy3kEa7vgb7fv6mFYYs7Za6nZ3mY4vq5sU9NL4VgEhu2YZSIUGdQt+qiWTAO
Erx/u7P1Tc5kSzYBNlqUbLZshvaPgNpBr/HEZIl9AiSX2uqnyogUOaTzvkJ5ZOvB
1A+QtgK2R2EVgMBT6WoK/5UGwbH9ldHNeJ9OTRV26m/cW5CaWnLJt3DfI1WIUaeR
2u+i22O+Tj5+AaMFUF06GSXyYC9rFKDX26V3Kr4FrtPIryYv/ddUjOpFCZLMBCtu
Jo68S6YpPSZF66BXKAuW0wA8qZVEDWBjpE5teQ9IPuR05WOt30/0xqTIEcgdDBL6
niSwuabukPendGyBOtld55KxxihocLSoRfZva2OgFBG3LXT2mBypbLE1Y/g8CK/c
PZq0Y+3TafJGNsHF6NBEnQBVLQ1HoJIFGFhiVa5oXSfuqOVG+vL3gMRsrnqOj0Ea
s+eHjOPcxau2Ovi6GJrE6EhucUK1sXkf/7YrBoW+R/YCdULxmddGjbycrzaUmP+x
EamxX9g5gxQwgvScoxvyantFnTFrXl4eUyuMvYMLfJ1hzjnyZS4F3W2w0kNpmd9f
2hAYxrcGCD29Qmk+7tP68l4zpUPB4QTCaI1RrynCPq5ue4rNjD5rlErPg1/HnZr9
ACheBTDMECfGtmM99wMFfkYbzGI9ePtrVcw05gbkBkVQkTbyFxv1P2gcf1ExygkO
OL611C4EQj9cyiDeNVbCwQ53Wo/fu3udqbO02UZFEXr4nxlbdbrZuRZYgxL8YjJR
oDMxleZDNu+gXNcl+wLzBXcuhu0txigAxFpu7NZekSAQPte9xDcZiCp4o4HorRNc
lOFXB2hlOuBL526ycNxlTGR5hPB+e6s/Ga1w1pQ93/KaLZBVPNIAX8jdgUnUBFNZ
nJY6NMoQ9f7xU31chSlSAo0EfXboFIr3VsZQnDd99RmFIAiswyjJSVXjcla4RX9U
QimJUO8sRVKUvcOYfBw1NDtvaZoeqg40Kn+FjGwo9t9lnJsl1zvxIDHTSyaYnGlI
+yn1bOgdlqbI30eM4oyq+TbM4HQh03XVh9Za1px0Ex7i6zNZJPwrTFuWf4xKXXYK
7IKWK4Wxplhgc7+9VQPccX35MssOnZ1cS3n0qo9GbyvKW4LfQ9URyR8nJseR4cRW
zpNuiun778VCEhNahfCQirWIKiX9YNPhhvugg3WlMxkv+o5jm3aa5uQe3bO2Tc78
tZSyvr9ItOvHNmN/+q2CcKagG20EaBjbLQY7MxtvJuqAR/XJMdmkH4pgQsdMvDlF
hW3JH7j4rVapflwxubl1xc2P7KR0ukV5TtsMlRKyoIMc3US7S+S4El/U9al5bSg/
bQRvONgef5zA2w08SIu+A09hAh2E2D9Lmad8Xl4qvJth8CWZztC78VDF1IRpHWMh
dx47S4CQAQ/21Hsq9JGI56zsPMR8s5vxOfrb1FQQmZMML1n1Drr7xtDry0gwPib4
DPErX0xuzkUytCGco+L6w18qBNFXQDvA9d9YEvPdTrXAdOOCaA66kKfVmKj1Oqdh
evhIhk9n6FiEVm26w89n431nkkncWW7L3w3WsDVtSkv/r5kHW+Fbv/LFpn6Mrar9
8DI7VChYndqbY59R41RtukX2vc0vTwSV0aMYAE0u7UwpSFhvxESwSKkmf6ePrXJI
qTy/gqUto18GTyYJXQd3ICiuWOesq3dnjjsK1Yj0t4mkdM/cZ+XR7gtVfI9gs3gr
/4f5e41VSjmPv2kOXJz7j4f75Lk4qaDO1rU9AcS+9atuozHMdhbtuceJPeE/61so
PTOftx/uGG5GjD96BPzYGnyg82gnJXmdSUervEFRtUZs3aku44jEWmtZJaRZ1R4K
wwbSPGk6Ghk9EKcaepWZWYA7amj3/Be2uciZlRdjHSwBoLVT4ua6T+drbQQmlnBY
t3TG0NtRr0x7TVMWZrKPYoLRT6YyJ4z39OmdccFUKxIjuZGPa0OUv6vhTMXGFxkO
SWxl4ul0IO5bkFJR4p7cXEhsEEzhKJP8ccuoIGs0DbPpUO0nxYI2AasxGNa/1yrx
jupSlEMaOR8/acoOq2qXzYEeonGYZshxVD5T0t+jjfP6AvMeG3JTqJivx6hCIPKa
v3TruzTfndfpCrXeDukcPfyre+A1GE+ZZTL7yBQiuZW7YQr1PRSdphQwLkHZ8ViC
jK6YmzoPa9mSaWV0rQ4p1pYMogAK9V8NJP7P2CKzgYdfSLJrffY9m4z/9VXHcUVB
vS9I0CGBiARoFIIvcJfTulJO0dXgq2PEzgDD8aysi5Gzvcy0CwMrDk2ftIyJLfi5
qNqtPSI88FvQx+46iKEXyVO2MB4NnAQ6J85txm1lCFLyIN5/SliDuufnUmb1VRW+
gd87I1459kf/GtbXyfiHVOkkC9a2gh3m9QDtNn8cmsc0mlUOkLS3MbKPYXuKTgNK
DoUkH/CT1VTpUHqysmS8FfcbJi3duwC8A8JZ7+U9xy+r0kAkeV0b7IlPDCuQo3aa
Q8DeInfxVyLba+QU7TUw5Nl7dhhKW34mNwOpCujtAGNU+CcgDosvwkShS4hyt+YZ
3hVGyePIZ4IOjE2h4XHDHjXzvo5Xh8NtAgqotAB6YFKq+uLXDjNpuD7+MRxPPYRT
mx7xQ+SlyQEiCykhvPq9QdSAOqVmS/eAWN3rWHIWLxTgQTtCQDePctZfeajM7dKK
1ChaIlm2w+abhhblRcfDg+RxW7l8vZAVF7ML88Wm0yFN80xKy5pX0Mi0RofpXU5G
WOIsdDvXqSw8fkZCsgscSMSD+ok4Hesq88s3+azx3jieIqqTRJ8hjMpWeOsdJd0I
Ub8UleRApioFG3xmv+9D0Q+ek/S9hAAyToAZcfD4BcEZN1F2IrUllRf5h+gGkt/3
JjcGUgwFQrseThDA9dMMk9bbiqK7Vuu7o/MQruz5nBGwjRPj0nTox+OmwgfF7zfZ
BQ8dyr7/CNf0vQWF0fmfyujuOp+RRUpQHYBh0QWrD99aTldJ6C1ixsIzU7997o2+
ujEGm4PS1I6JiZj+jwpx2acPORMTDio/GoUEZ+z3gXzKv8oQJOwK00gu2xWsHJXv
9VjnKqQBzxLaJF9o1q1EOZRMs83Nd8w9m2POs9wOdP8matXlIyJKh5uov9vDsOUb
Gffd9R8hJNRUnedRMS81YO1DviB1ft4GZt4jGAAhou3M9GpYMhHx2hZilM8AK6hC
JMUvTbsXZEzwDkCKoz9uNI4wkpVEedIH4jS+TsBYT5sM/U7qfkq7TIoEsrKwtis5
MbzYTAWkqInnLKueXNrWvfeNFMCF7rd46E/Y2g33hnHTNR5yo3LLZmpihVT5A7jh
tjekzTIWIWmaRPOiA7c+0QWu9KsIQqB9Lcvv6S31jKzlakV0m949sTlBpzvGWm9G
RX/ZmeiDYhqC+uivYIXpiK+RJmvjFZnCWIqhDIo66x2RmFxcfw8l2jWkQc+mDOpE
a+0jeqMFgQD1xVsUb+9rkgh4d5Bn1d3pPjXYSl6ZWKAHXahkZomcwyvC60MMvfZD
L6DyhrZIvZwg7pDtbytcxXCt5Vl4wedUisEan4MdZgRZdVzztErcDyce3Sg/qlHS
J37/ufw3oRKY2QdGek8VHEteJRnQ4sIPYKx3zhWSR981qn8fHC9fOSYrqcvbPiM9
kYmxW8SpkXMR5nLaRruFchLVmUGPapdGJT8O6bGUBkvhaSW/e6MAlPJ282P5VKBd
5gIL/8HDu0t209ErZ2rcNO/N3rVgzBolzOqA18Yw8RgHGXQyZL5mSNmyv7t170XW
Vj9pi784nRD87DWxRtnHLlt9YYbNINR4q6s5p0v9EcEM3S+YhRpMZkMaiblpaQzj
QaijCXew7VGqHniXrlx6XGHjPwcuRNprOOETszgksOSr6Gon1sv67Rita6Tlxdx1
sK5tTuHoqhBBQ7pDKE98QqqyFhjnaNH3KgIOeDz6H4wlxLuGZv0R6p+ZPr4cMTxm
vhpAyiOGeXVNU+I1yI+bjetyAAqaqgxS7a4NRuQuBDz6Q94BVbL3GK0WcoEtxJVs
XC/BnXlYByNwbuhh4a8upmpmQ+2AALexaGbShF8da96cK2VRcR9Eu/OqtRfRQ6eD
74QOqhjGjtcJqZrI/VzxsvXzD+8WCL0URFbd97XVDbISWTWPReUKFOLe+2i9RIfg
auXMaN6jfPTefbFbCKW/lbnrdTUFv+t2rfH9kF6QSrLqkwZ9I5SfYpzBfv/UKOVw
X4vZ5etH6dkQOmvtZYcb661R95tNG/nHmqHFee4ltFA1deyjsPuWT6fcyPa6LyA5
WBXKKLifcaSedtydrH3YqSnDlLsl3czg+QxnG+OYPEgb/Na5i2z0BQOQ5r34rJU9
R0xmQra36MbCvZQqn0o2X/lkzRuYXaXp42otYN7YdelV7dwpdjgGanl7byUaikJq
eCLP0iftMyX6BywSS1EJAaUfVcHsEbZDkIoZNiQvs31tlKjpRD8/gyLXEnDgggTx
3uK4bWL++DwV3+WOhvFfD01ziZRfvn37P6P7zduIRyh7xico7H/9xKnyVv7vFVws
N7jpd7rjdvI+FnMmbPMO9OIlmGPBht71nW8M2smzwD5avAw6JeSK3OVMOKEEFzSF
qN4dRVpA6otNsaxWxQCD2AkQPoA4//lfJHhOHRM/KetmtQe555PWJI8kJGXU8Ll2
G5Eaa9HucHT88aIhPdqtP3a2T+s/QXjBf9qTu3Cu0/ANRZFKsDFUZMCdF3Wlqw36
LextKKBABbeQJXOQyO5VLmR2qQ1MZiCyV3uO3dGPL4GMfN7C7F/tumyp3epPAHO9
nmERp3exdaBNyaUDrDq9+iR33uLxXHiv046v3CsH0Y7bZmEf1QsgnTr6/NjMMnrf
Ueoejx08MRRAmP23o4KgSdzn1MQJcGolyOShwBkS94A5DeDc5mUytqXeA9bwOPq/
vVNV/AG/IMdP2G7lejyHZW3wKUybX2YRu/NuJwSGpFTJGmdAFSc7m8RV38LAqjwv
RyA7e6Ggelq9qhFN8IGP6vBxugK9AS+wteX/NG8FUWwJ7A0SnMJE+fm7Tgv2WKBK
PmqNZw/1g54GtW9otLO1g5PI5jG1831JtyeRTIns860a9mN1QW9gAkwfV3upsVHk
kOGAOC9I6tv6JrAh02GUMwh+VH3CrVOm4joA5dZPJ/H2izGuvy8QsUeo58TBTb0J
OtpYmaoaKyhWoVZ+S+81rqtfFaHQoMTTak2fjiuAFkk8yxlRZOe8W7tfXvymCPfP
g1x2MrA2AFICNBi/B5pf0020SmtI1BcuZ7aJxS7WeL4UbJPd4haoVPRccGq2TakW
AJPqx1CCPt1ieA0sUcMWMV5MrgARhOtXC6cRBaT8J5xzyJZKP14AMPawsxi6dTeY
laTinGKfGpSfyxMHU4Iy8qzykQCHlKhj8uwLsdQWvXnXriPTT5D936Oa9i79Iz0P
QbgwAfoQMkkvA+y85xTibkolRF8zxRzTNVpKDTRrlxO1n8X3MLr/qPI5v9JstVe+
irWMLI7Ldiu50fHjhBZeyWsi8MKeELofJzOZV3Uefq++dT1rmzLfiK0MU0aOBKbE
fZRyKqF5wbziDsGI9PU42nVhLrRbPBgvKkAAPkFWBIch6yvE+VwrULlPtM6AExy8
F2zvoENXgCM7Avz9zWPqrmOCA50e6+sWE3LcX48Tx+zDMTfbc87I1cVQpxQ5B6kW
IigQdn/iVFhjCdO2veVcmQrzaZLHcY4oaZUl5KkYLTSNy2qgNy4DFMiX4m3mEj5P
4qJ5pVXL0xnoK4+eMJfB3mHJtrxw61L//6Y0bL4dY+9PhOxe8MnAr6jmxj5BXc1r
s+weZ3ARMhZirbhYwRxna46Usm8kIp3X0PvJpeXVB4CfVnWTxMA64jqg3tcPiFsV
cP/7xvVlPQbLJqY5Zbpebv6jAM5zsBclO/sfyOn8gjjzMBB64vx9C36me0gA2UN0
nExvoQ9QDLw+JnnWx/5HQUUgGcLYH0909QEMef44c+ue0uCAZ2p64gdfO6JZeCBN
K5MsZM17NM4v6FPnSYB8sEr2+F5BNkSKyTFPdKWO1fTwvc2I42GZKbN7vyMVq5zN
+8V3P2L9VlPXMZO7GzW6kBL250a3um2V8H2aqc5+7tY0P4X0T+hMxje7fJQwqAfX
ceeJBcv/4+mihTGUcMMqWlh6LDR6T79rfFSCoiF4SW3BNs32wz8mzwsIng3lCCAE
V7u4SBY8JfbkuStSYZ6kku0jTX0qJSoHNShwuily+wbB4tyZbLk2Q43MKD35/5Tn
Pa4tg2ef7hK1awf0gwCgipMsuDVfnUZv1Mrji1Q6waJih0JlvWPTRxw1LP4XeDF5
iTV3GL97nHp26inUwWoaV1uQ9da4uMZGvcJXh2x7KyrL4OEZu+qU5TSyBCD31ZoK
89OrNEMycjFO4L+ttzObctzMG24MXe9FlmWgHC1jW8uYI05SH/bGoIRBMvWH/yXg
bx632mxTB3ibl9cdn6BtUqBVeVyPZHlwrlok4X/Odt4gnN4157KXI1b5t1gvIj3V
YgFeaO7oB07HZBkgmkgf6qQXqSj5ttwjqYwtOztNWjUuFGRGAN9zaVJNQMcC/WzY
ZkE40a46D8KGekq6OtmMqh8w3ALa6nmg0C0aDd2OKvL4kR0MSLluteB2HNDwJW7P
bJWwV83GegnqOMeLOILetqViheTEvlRgEvVojRwJfvZRpcpW4OjCz04ehUJd6m6l
XLkimvWrjvXt2DLGBvm5xSazMEGfyTfGLoiKc7ay67ebnbHDzQ8NwyLfHuQS293c
8Twadeco38GZHhGmqRmrBSGmtRLVZAi1SflT3toeTR7JSAUZj1mM7xvFggWYM1gR
PwTkF5GnN+/grb7C85LyDu3niXthty92ha73QVkDaZZt/bbA+KlifZTHiN6LFEpp
XlpITGfX9RgTZoOvDJ6yUMEwgzuFhD2nhHLJ800CT5rkZ0e8ZQBh/5jdtBsiyX+q
GKwTnY/Ta6tzT9wxBMnkPxM12c/BOH9p10sntob9lwNrclmo13xqbESgVPqLUfdX
89kYuX6xgKAmjNGUlp1ts85VSDqFm+wcHoujV+GLAjz500tMUXarEZ0nOHzacEtj
L+CQboadw/k7MZAbtyvVLwTJEQOwbnABI9H0GxK0dLN9kyuAPsafiyME1PeGOSpX
c0gnZZQ8XVpwHivnP+K2jZal+2PEgpYy+FobOLvAt6qRNLbQmI4i8gNPOOeNf2Qq
eSbB81hUwgzo526i4ZJsZhSk0rTNdk3ebh36S9pEGFaf1aeGZgvE6RL629S+DctL
yJ/7eKH/ebv4q4fKBeRMCRKrWmFxLSs4RukmWB9gxn2xizO9iEkt9RsCWVypk7vq
oUjXOl74dcj/aWv8/wwczgSVHI2DXmIMccYdT8NS/UGjsRPD0OFVXk4wuhCI88XW
s2moBx+ZYWZiJhTgxI/kg4FsUl6g3vEsO6j1JQZOCsJH7SP4pAQB40WbBmye5Mgg
AlLLKqyh/GROijesIsq0Xy7ahQ5ZVOQlPh74wMreG6orM7a288JsiosM+RtLRxEO
c1c4oCtzlhPceUadGhz7K408Vl8SN4BbwCG8z1UAEHczspUyqIVx/4K9/IoQsNNU
1Px7irVg1Jl9nu0j7JSBUgoLTWj1HuAUvGnJhhHcSJ8ihSdFJlMcenM05cAE46mA
eZTtXCLvBiLBzdI8ra06nk/fiE8kmqVM3Bz6S8CrvvqUKKnzS+fKiIKcLDDgntHz
7XPtOdPjkNJJ1jn4oQeZKs5DipL1C9+Ro47FmMfcEGK5ihy+pyvDzyQwpNX+tsJk
L57yxw1Dn51DRNRcnyyN19M/GUc8cZg4iajeeCRahCosI/b4nqRMQ2+5OttTciap
f4oxQ9/CP9eZe4HqVwZvGJhf5TYlUBeyXaPeuLEqoF6WgfxTfeVXy1VizMiT0bNF
VxdQzniYyPEhOKuM3ex6AKJhrAQFxXYVTw9QO3hH+6YpmoricyFXCiEFKFV4RUSq
ys34c9RbnxsNgycw41nqaS3lSQUvh0+M1RJ13oF6AfT5eolnTz6jsiEJGfmyl6g5
ZQheUIpLgkRLAfVUBYQXB469g6w7poUV23CUgfdaJ6iAQRSKBMwXEFhUUBkFsuqt
FjhWvPqT/IUnR1ik/CXJJdXqi/cNhxYZYWt7q638/33viaWOFid8StS9cg55J78W
bLE5x2xi0fbd/M2FrLKyPF4wAg+2q0sKVgtyKJSoY7u4RKm9kHspC+JJwTVTu12I
IH9IZJ2AKwBMisOp7HBGM1S7gRAOq4FZ9TRZyCFuP9kZ3hNJ5xgjTY3guz+WeTHK
20eRVOOBRZoyNVUOsmqQcfvV/z73fS1tbL9d1lDIEcEJ9dKFxrZqISDLqKBJrHtj
PyFrhX4dchPKPkZv0pS1JtQRpSZrg5U9t32vKpG/BrB2Lh+DDHQLy/1HaOC4X7Ry
46rC90rTgHnDjYekNDWkSrMn3MzAlnU0fUxXTq9vTGJ8RLXrHI2L2iDC34jGsbdi
ETShAbgAUrZtLg6zwoh1+VPoQaOhtIDkqplIG1ZFoG0VDCi3rNG1hu/nceARrTlI
tOYd/XyYkQcT5D3OuqktUgM7zuh9l0t14i8aHdderwziP4I3xn3eJaLBHfka/wU9
M17Kivlzvq4SnGcWyftZiEoR6tKsd5o6IUasMcdNtJ+qhBbp8NuMSmMw8he4Zmjk
pIoxovJ3z3doF4+HPu1HAMDWoMUXuaZaMZDUFGjer0iuP9z3SazG0TFvTlo7amLH
0f48SavZsJWsSnJC70PahUONur8yFr+DBMJBbNduH31Z+VI7zJCWEq8+1RbCI+nT
jbSeov75mWgIE3bzVqD6XvF+poAewmckSoe62shIKbiYH/YPP0sZUSIbItbYs9AV
tZfGjPOkB4Ir5KHsaOk8SsWCsoP/RHQBEwgmDQ63RvP4S89N1L3qIKtm628gv9pP
d/I2CXCYlhdh5r/XCA6YRqq3m0HFZH9eOLYqAiYiC+Hp7mEe5xGYHiu2gTKpgbXC
E0r14Db/FK23CcsspiLqgCY0bj/NE8uyE245Lm3tQWPytlKSradRV6YRIiTvOZFH
/jCu72y2mdR8ywcixEOZxg/NybVNPPw0TGQBH1k3gnoCrVS7j3WbU9iFWc23n0Vi
EXAg/iZ37NKlWs0Cx9VIoS7WE6edrz4Lo47Rhr1QNpc6sVLqiHJslEFTmHFih/+z
CY8ev+kEv8sr3CqjHb4Xs5BWdU6l9sALt0IcaKBslVWimqFscwSfAXLtNkZPe8XC
7CoKdH4tY16HjzwsjsVAyh4jH1OJ5i8Ua2FQVeQpZBQq450ssilbndSsrnvX2dZx
bun1JnFpaXjVq0zfZ50ZuuyKydUk/n1PjFTGEPWd12QBfO2EjxRs9+J0zwT3ygE0
AqmSCry/vfJDGRXJ/LAvrGWl2/GypfVg/DXmGYCa6VvHC8+4kvRJ0YYtiM2LtvkX
sXmWunDD6/hJLFx3WPo5eWf9Bo4cws0531ZX2iEyrpvy7ageIE1qFjYE0SDL0+tF
DJnDIamyK+yTvBlRAbDlNem+N7rd70TBuSQE6WvYRpyoCGy0Avre0sdKk60jlYnQ
KhdgswVSobwf2a1WwRwdA4/AVQvytqpGgLe18/DYa92UWdeFOq77LFuqWu3g29Rj
wlyDPcR3LTUw/Pws+lNUFBodIz2Jq6ALD6FfvOSHG7hNF21K0DjSBJza+0Mcfw/+
8me2KlTDJX55VWQnKvtUypkYHeWbLLuSMoceBJ/TVaX2KjhJ34ZH9P5piEgPHOx5
89t5JZYTqsf8eXO7OD5f2W10HC3lrj8Ed3xloXlS7BAzZrgOSFqnzF4E20m6kky0
MEunK7fr0RmDvBSX89yU/hIgwF7dohe/JSSi0yU4/JBJcOJ2UYgqfLDbDLThvzpc
Z6tf3On0HrRpITR2ofa5WR7UOAODW3nRugs7i8wMsiEgIW0juZnVFcnOwH9ZfAaW
o530qc36ztbJv5ionnZn9GK7LXMvpgJHOakQHWwzu5TQjdyjYrx1VukrlYF9RbmR
mUR7AneJ1iiqPhm4DFq44PK+eWSm1yzZrBOh2jCHQjWlR08xx1nl8MW5CaAfgN44
jKS6UwE8FIF1tuDGIfHUzvH3Dofqp8/Z/Cd1YQOn8WUezmcRrvsdyfMqGPTzhs1H
AnCT2drNJxh96p9LUYGC9FNqsxVTH4Pr4KTw2FFTPOkCFgr6t9DWX778BvW/qwMC
uX/2/U4+S5+BiMvH1D0gANjc3V4XTm2u9oJoGySJ+zFmm2He1ZLP+ATzQizqXMkj
dOSe8rJRUXd1wNEFoA/iT4zSOAD4951Wcxz0e7D2vGQgeZZLZ0rGNy5QCen+VEpI
m23FmkSMYUFy3/0EKkt/0z5fXtYbIS61GhlOQa/6gop9L5BKJOWaY9KRfQNF3BDY
3i8dwUKW6LFnwBlyvpwa0TZXjhqXOt94tr+QVBjCTgyGEmuPpsJr4Q+m7E5XuMHm
WpCPSAAqycX3AHepUP5YmUEOzQT8ZxPKOdihqrb16D1PqhTkA5zBPN0x2dv9lCK+
sYi8V8wH2SrU4UnOPMVGz0XJ4VdCQPXeBF0rw+UCpBvYtwD6416AyKKfws+Gy6GD
UL4iMfBV+Ue1uNt6vwl9QEAGGlUiPkVSMlI5uPO4tqwQrLnb6piOceWUdQix0r4F
jbzJesQIoZ0oHEEVujHMluoeatNw+2d4vQTb8iOrk/Cp3I1ShwTTw+5Hqx2OzO1B
wNVJOoMMvkCwj78ek0CJO8Tt9UJDlTmBhiP2UeNt1URy0QcGSy6GS5PlYKfJsRp1
bVeTohZYA46PMvJmzi48X/UAxcLUQN2LYDXkara5JK0vNEhN5TA6S3f39zrIQx1c
RwOFFy5a/OnX8j1CelG8zjqNzsDByG4sVsqA/iDNz/ZscYNph5rkT3jiQSYRDyEn
v8ym/dp/ZlspcWjGurO/8B1UtIuTePs67mr+l3QEuFNcOwif+juTlCgEKJLVOlD4
GmzCV++9C7QqWNW6eYIemHjvgktevQBK9uc1iyP0GxoHuReJculq9GcPvmVkyeDp
2i24oW16t+qJAryO0qfLaeRrpUMx+XkrwFiUFAyKgfs3Hs74NVbYgP/SKwQN71aA
ywFyqELQ/iV3DEahpUnwnX2yi1+9IVa5VEs9DqiJAIWygBqm7J2COZ36h0y80SCR
lWAIJyQG7E/8+ah5YpKdQZr+InvqxTXZ66eliyxWZBwvwbnnn8LJTfTJoCLwq0T6
zbJoJGKpIvLIVvwBI9n5/mUhqriGaPrLVUxQof2PaIh2rxskWF0zHjE7hllYCy6b
/bhSX7vlnstzIwPBhm0dceTuJgeWvGGzceruCtstKxAjEiWo7f24LgqtK7KhnavE
m+ubM+pnfZTOmAK6tujJDVRNTDKaJhvQdfGDbhawpSp/JRtll3vM8z+gFT/m4zAT
ciZpI/XBBl79+4YoSfKS60IQVBZsmYijPMa1F0S2nVjnorQKXAnutxUVyfHNCZoc
Dyb6FjnDRZzLXr2AWZaH1PXA28aWAyOwdi34qQDxR+vpvjThERlPMeeiIaFLUPld
F4CjzJe8uqenllyOpsMWqDJoSXHq060uh6I9Fz2rb/8nLBtbZVm86aO0BXp/nR2c
Kf62M4fFBTpeiXp9nRzZttJaQs4SGnZYABWW7ujSa2luzMgSdMZEI7+xAcikXjCb
7UHRX7KpA4xwFgCWtNGbP6Q4sPXrhvZ7Ob4R535jUnUmcyhzMF3RQdMHu0zD5nA8
cLUXci8T7Jo0orRyw/t7QVn3vFbSghG/GYQvsdPwGHK7t1en2RCXTcz/EVDQMfPY
tGoaDBbJRVEbDSDx3/f0pEMYj8uGOTwTSeezP0NeMfBeS1C+URP8V8d+tsP4h/yf
eJuL9KTopmaYeKIoFSe2Ve0Eu31EwdV9UtwkznhCKJMPDq45q4lUqrgIKy9CmMOn
RPPf4YSj7u+zQL57pEqMJdZmLMmfCTeRbJuuzu1bqMYj+mlWOPkROWSee6yA8Tx4
O9/M9DPqtzbNK1iSsN1a+y4p4uqzXDfp82enJPR9zVYTzuVRnGqG5o2wtieLSBot
Zidp5UWyIgnZyMu3KXPKcmeVX4hlxl4AhfcQjvoZYYK7EP07KYmvRNiX9NuIOVF0
Hu9ON099ldZNels+I0oKdXDZ79+VAjpSL+kZ7MOMpi7Lpcp3/73wBn2f9WQIVlPi
FVM+kXipzhPsVGGG1VLf5YJk/xODNeRsTtyQAGD59yEBpXFi8XdM1vYdJOBueP7o
rsysTaT5PIzu5mTc0PNeWD+D9FGw449RC2XjiqZ0YA+Y9JUIqvqJdVNmfXhoZgtW
FTF4R/VoBhUB8nuzVKr+GOkSmkmqJB3o2KGPtMwBrnGEWtvx5Eff61GsyC9lRV07
quMHq3M0iSRr/+Q86usBeYMpLAuA+c6Y0gk6y/d51VFBNJmLULlBkrlqQ2Ar2gWD
ZtVIdl87wKYF3kQr7Xlpoq+crRWI08flMgr0SAj6xO6bZE3+7u8cQjWeojMs2DWm
V9WeeSCCm4ZVvjGyfV4fLHJTFVDZNHJrKsRO34rqtmOfDaKSlVCDZd5QGuWqhKl2
kiAtTPJ31IgfrKUQdAqxpTojC40uOWSLJ6V67uaen2zVBbPt0pPZQjojHAs3aICO
oIZmIB0SzoCubOdIrAOb18bRX4+OttVPDAfxlBTEHgO6uSwJaq9Iefz33NgAOI80
4dkHYJWTY47qVbGmhxJwiSnGHBWh1D7ZzfkaB8+85aFpIhpTgenqrTu9RG44+zAF
tm8TdNM4Xtkh1w4GfI+7hwglovOeQ1Vp9q6uWtnze5nniJ0OTxclnSvLD2QCAUDv
LQVAO+ur1C2kQvWdNuBfWmUxWvol/iYkehmhkhJv0AewV0GJU9OR34j9Hbw0J8PV
o1XiXoxR5/LobnTdXNOQCBuSM4c6eu7JAmfrGHDvtnBydwukrWpxEDWwZozOt/ts
qXpS6XVR5Zf/eoVDLmsHimvoO4d1yxTf2pyx45wwXyF2k3mR/Eq0FVVLe5WmJvuE
U21DASuv7dZcLP1zRHsniC+taI26M/2PnW/2yq0tFyw7N5BEU3JOBK8mpV2lID9b
Dm86xqB2de93kDkM6G2TKIMYkxSwQ1iwXx2K/ZmxvdwJOsnSw9j/APCI+C7ZVsPr
G+O/Vfh3Zrrzt5FamxdB8B16XK5ZYeLDRHX22lm05P5glSkS9GhZaOnp7Quz7UIc
E16V4MTZDMqi/aW2l7osgVgcMe4KHzDcAM6PP63dKA+uo9PXxxcmjFLR8TIO0IWm
a5q1a/z338AH4kvpeh8fkWr36LLkQJPWesLtRdzPp14RPfwcDOCMeI0Upkf3qDVK
V2fD7cQgds7Mgki1PeRf4bbb2JlOqX2b2FmUhIc+MQXst+iL55l5WlvAluvENbI1
RXP/ZqU/NSe3G7t4nn2NrDN1OCq+/0d2pGClutRU/BQoMuf296ToaXNC+xXzuk6l
VIqL2sJE/+8DZ+mfF+KuJ3Fer46DdEVzR+3xz80x3EhRG6wGEokrlscu+UvTp7kr
Rpbp2gs1zidZwixnd2pHMIJYr25pOl1WVdNsZtmktrE8mQp5yqZ84Uir1XvCBO4j
L/x/7M56Khifc8JoG2+n9bd3pq9OhFzoepkiU3HasrQGIVQ5qSXm9Xg9oeUUMtFQ
JTVDNVItMUEXGCjMiXXqlMNhet1Uqn9yhxdca7QnFoi32Cey7QZoDzLG0c1YETEq
cFQjrT4wUUqAAUu+t6x+RSx76zwVrK7k19GcCh/Qz2zGI/pIBlQY5ERoxEe2HPYg
ZGYWQMVSdloERUxxi4DXkZAS653sQvCMHApSDrMbRBz3uWeRKYBPOnAYVBJF6e0L
i+Ntj4rrly1bl+m52xGhEm92Y7Weyo7ZcfbYmIhBQeUNTH3YXSi73PsKm0J706Xj
uFEA+7geI8KTV5R3GisngOoY66+ZzFUbpc2xE6yip4e+JD7m6pYJTegQc9IdcYMo
qzmyeD2PpgtFzFMhkPNcZs5jyroXVR9g5/R4591GPMosbccD/avFAmdUdIY1jjWs
X9uDqkipwaCuHEmvhaeRwNrq6lK80otuU4KYFpv18pjxQ4Bn32f/llG44qbAc+FB
k02Vvl+8bU6Qhl4BxuKkoIuv/rDSOONzQk+G4taSyfGWQ1qzyelODchdbjtQpunS
7W5Gb76721Q5GUKlj+LW4eKBN25Acg7t+CvMM9uizRcN2NrrxuuyBjm5/FrvBuRs
60Z+5oTdLpBRL4IRrzhQVoR+bFR0ZGXlYbWkBzB4gENfKhiMIzxvsF3J/WOH649a
60uAfnNnlRG8pB5zNLa4W1dLo2csMqhUqer8qL9C/sS/ych/ux+gRpJ4pPHPdP1W
Lv1BVEreZW+eNKF3Re1MyRPhVJu1p7CIw2RTFpicoPAX8lZAaUSGpdeU9J5RPXHo
HTqrlJeDQXCKpYn8E+RoJjIF+biSui7Dvrr3VItsmcxWDhkDpWdJ5nCX8wAV242j
yIm0ALjjT4+LFkMRnphEDLynQZsQ3JJsuRaRaSXJZTWZIV/mRKRqXrM+SnpOH7ld
eO5OzzP1IdISxC/+yNZa61XYhbfdJ+QEHGySURGrm/UlMYDZJIk9wNaXb8PTmQS4
dbC8KePzz/FHxC/bKZZpR1PBJ5uYsS4SI4LY0TzAPtWsTIDnMKkl+2KbqH5iYpLH
N5UjFcVdDXVRRhJuHPfWnAQgj6463ewNpNr3at1Rij8xXWjAzu8hNUAHNT+vZcMj
NX7GB0c3wNurxm/kDNCWMrSa9FCMJNowQdUKCY6NTGt7o5fMm+jjGL7lgIGbWYDE
OqrkAc1+5+WZ9dFwng+hWdVNvzBnXVoDJPQpxqnMgBXY4nKYIpAh1GkxMww5GbJT
nBvS8TY+DeKTRJ0ISTKZ8RBx7ks4XNHE1T+Plb8g/es2VCbNe4nrkDxiuLN7SrgM
QGgP4Ecx+ufpiHVazcTIIC/4Gxpb0R3Mmvnsp0ISd24lmKcV4oBn9sLzDYAXiitP
/5efSPIioNZNbmexUkpXfBRoz7o3UYV2NI59boQtx9sKO4wZgSuHnhNu007WhqWB
t/HV0rF0s4fENER937fiLNClwI9yrP/qHO8r0G6042Fhb/gsa3vNYaq7BHMw2+1+
TjUSYqtlp8AYdQvi5uC0YWvlwm2UONxbgeYLqLvbr5nZen5teiuG4AKrT9KFdlSB
77eUSkyEzuLRsjCaENAyus/vg53N5Vo49c1xsnolfm2batRsATKvmXh+rCS2cNN0
JqptCiX7Jf4m8hXosXJS8FD13G8z0LuCU0mscN3o5i5Qh2ch+VAQiMqoDxttit3l
uS/jB4D386CJyBPxYM4XW+q83YoK6VvyNrcuQcpsK6mcexNNccbtpx2WVz1nK9tB
sUYmWVUjo22ai376JbuIV1DskBwC5jAHq6rDb+64w0mxeqwLOcVzTen6XLyK5Yg5
0TkmOnjfVxvuzm6peNWkoH4FbfpLCdsUywpZjF2GFSzGrslKv68eW5RVGInDf78n
afBjjvRl0cM1ZgJ/IvtLhR2XdGjo5U2MkFELjHOJg/eKkt61z53ShOTxuZmWGFD3
eMI75BCt1MiJ8e4kvw82peMGB10cAHwoAQNmAOF6R4AvGLoQ0F0M4Dbt4nN09vcB
xRzSwoD052/XvxyHO2ZV5ptmExE+cWAGOG0odCca7RIYiEFicL3JBoJpjMFqevuw
nP/DpvZn6LdcHiMbHAtBgunKZbH8D4tm7U5eLsC8Eiy/iF2T2Aze9+/we/ixjgKD
+FB2p+lb2OEAxgJyVE67wfvvcqewSlW/V4eMmpbxqK0hn9VS37R5vOlolf6hL7kD
Kdm4XcOIAkMqMM11fo7ra2TYK16I+r8qYRigy0F/PTY4ltcAdNiMQMVAdekmX1J0
rL15ZH3sFtdwfmADU+lt6rFWmt2wvKKA297SospAMkXbRlnKev+wTN4nieS4msNB
kZx2BlsaXzEUqqQotvwv2l2pLQ/pBSc217hV8erhXxIixDMCX6XTYlW6uOLTOjaz
/vO77EX5i6ABqGMB+cLSCA614dww+cWDldCnz6rpxulw/aaOxXhe5+V8GKJved6m
ywcfFbtYC+8Htxbu7QJbDTSi5gbLZNfWVH/1/FPSBXMUA57KG6pLyZsMrRrw8+u0
q88m4qz6BA2cIqY54BAuN/WwYuKNiTOOW19x4aw2kzidraYqH5AOuXGdgZu9M9vp
46r6h+OyVpiTW6pACAf2Jp1noPiY48UeeyaCSn5i2UfGrZqBtSf5YThGX80xwI51
Aay3DLgWAm1Jx9ZsDi1FOErp3hM215ckEu0GyGE4+0IC327w1FUYkbewAbRBuOn3
Dg9+82QS9s7JWotDLChEh0qiXo5YyaniPuhDg+MUaia98ebNaXCHFehOfII89fQL
03yS+YWDjokyj2nol2pQhJX5iiBiB6p2UkAZlHZEb/uECQ/JGd94nyDd8SsdOxJ2
0mu63TFRSzTi/lekbgIPlvmhYlfsU7+FsOHUEMpXU3wrQCWztlx5m5cByE2L2Y2U
6XvflJTL1sEq530NbDPuKqKyCbht/manmtiVSQaGZ49QHR45nbWaBE+43nJIIAra
4q1g5xHTjPsTFyBBtx0uLLdBCLwZHmCBl7r5LMGxf0cLazpeGxesyx2ZmMlKERo1
BxfGd/D5X6+9xFs4nIHA8Rb9LY2sTJFCloxeNSJlZyX1maYSdEflYC/o/JGiSxa1
rZzbEZXbJLItBl5wE5s+4c+mxTecGnXNAZq4+QBPA4q4rYLXXhDaFNx/83gkbnxT
qSAP+GbmMFrL+qmexEzHtoMd0+XATiCCV2aYeeTv2HPRRYwJnXbQdjdxCILN5OZo
4sAa5Gu3Y6SgmZJCl/vyD3kL46rXSAmc5tygeGNXxEZmzbScIM+0KQAiQHcqLe0+
Gxwg/Wx/z79I/767dw4MnJLoEQg/jt6nlpBrAdWkboUhbdMS9YwgMpUCoaH8OZTo
fLcz1zXD4vFA4IRfh93tEmFKwP04zt26VH9A1WaNxPQtlhASudSDFKK1n5n39ja+
mFxW1M5haMORzgz+n/+tXcd9MCWOpOxe7tryZVT1Znw6dn4ukb6TgsHJOuWv8mcD
6xQa8O2Pv0xXaCgodR2QR2o9v3QT1No87iKksm7ykpU/3b8NVDEjwPXKHuXhekK0
DNelWd9q57aAO2yG7NcstBsBPpFufH/DWIK+HzjXnuQfEUTaEoMjSaK27gtXmbPL
tRSQlFwZdugX9WGAWXEthFDQRrgHjikwxMFjfm+UktAsRU1sxKIXg45/UZXvOkqp
j2MuDohaDh2u325Dc/A3EvkUOOWd6RN88+kyZoDNB128gkZjahUaM+Iu7llpRCN0
hHlaIg0kY4GyKNvfIBq0k540OlDE3XzLexLUk6lw0ajXlMM8bqozzX9G92Xex8Sp
jzKCr3jrYBYn2IuKuII//5ypRlfytGMQPyf5CN8bMgsVWfQTrw3x0MrHl/3GrVIG
PLUKZkuzB+Upx7+jnQjLKp6qhUvkM0fYrEP/KYQ0tugGdoMrnoR8iwlHhd46mcan
Q74sxphUVhFtSn01xNRmqGCC5X4EcdFtbpK5um4UzZ3c4P3tOEF6IXcfIw6TLwVR
DWiU2/LwrgiiwiT+n9Z+Y/4VnNQ204EAlfgG/Jy0ur0IXHBVuodDC8pi604xl4iY
lbvM1l89920uZlImvyCLheN2M+dUdeMolWYIAFI3lPYQbLrcNGSm7NWMit4/7Soy
G/gIfjkueDnrip+qp3ewgsc9Xu9fyLNSaCsrYCIe/M78jg8KEaEgzeMrtSL1qnid
8235BX7IgwFt3sLRaNXaRIYZdTL38Gh04yiQ4MHPkPhMrrFDKgLWNV4TD/IA+KjT
kmxWUoqGHfNk78zawnY95fsPUELteR7sNGjGf4ryL8m3UrO0uwtFRoTm46B+b4er
MGoLPjbKMdDo2hBcZ9+kenwwH65sve9+fzGtVtP3RqqJlM6wL9M/9PP9qzCI0oBX
ro1fo4njltnazdsHXPvAyDsHN/0Dxm2uLXSpzy2uxaa6yzRF9+x5zyPisHO4fC51
na46tyKmCaGnFqFmxXkfbcFALtgBXAwUnfS7i4oTTjFVQMoOkzjR5nBJLonxFbWe
hK3qQyawCpy+C2VyY5doET7Bqc5jz804XEUowzb7QjSX/Wo/x1YQZXpRE4P/kGBH
DejTlcVlDlZD6NLXz3NtZaFJE9f4NnXDG0j6gG4KU01aIjnuJqf3ZI3X7DSNhR+I
whhIaj7eARsZRaZnJ0vtjAVloX7K1VwPY+toq22g9+WU6SNjx/8UfZmOFWmeKXsB
SRnFM203nctC4OaJLuCIR5n1+WtWuCsGCglyEj9AGfQczPsez8h8Hhcwg7uajqaZ
vWMgf090CsyWEFb4reJqn6ekuDHkB8WzMFfWD329eXI2nyoZqP2HSpQ933qA8lXz
vNi2mZbFkgbSW4Ryz+qZQUrEH7GRtPiQqIo+paqqI8cS0k1uxi0hQH6kqDmETIgB
3hjd3kUl6lLOXUD7IhwqUDhphk4EYwl6Zn1yGFN11DtuHjT07VVVVhuILOhV68wC
AAtOBIzkDO+FXXi26qL8YdLhzfS18JXD2nTZnfKUCxyZfZrXE83Y0Bi+Ha3fvUo0
w1VQRNUClm1b+yj3NBIbbmxVH2HyeFwUWaJVrwKtgJzlkBE5fZSapKGDkH/CmriU
NnG2KnxeFnbSzu7Tq8Le1vzdkArWWfF4wFf+4Y74gf93M45jEqSAjSP5av2JThNy
1ZJz0SgNxX979R7A/Zf6Wvc4QBQHyfYmMftPcUcnJVqsuYVPPRJkN3si2zeV/3Fg
PRVil6nANnggYsI5FZ2ThbS7xxqgDG4xYUHj20EpAwhtnzwmPyT6ocSVqeAJE5/Q
6db+xmat979z8pMPaHc9c4OXZFI08YN/ap3AxZxPxhi7gV9CmWtBZc+EMgsO7sIs
AOzgp0Khn39H0nUMt7+P7ruTAZ1m4Qx8ZYhahP8Q819tfN9Rxy9MsZxtpIAiGStQ
nKRU/W23oQahxjSz625wz3jut2FBscOIBXCna8l1Wq3VrdxTeKxgEtrZkQEBRl1a
FbnzFSRmDpkby1q29yEmX0GPES6g/fmKp2CmmsVr8CEkCqnvoUmt0Y60hFFrDsJ9
TmjyqI8GIA5qy654ZJaYI65MKwzLz9HuB4K8xgmajnlIvHgVdbUaPgUTqWb77Po/
xiZUvbOSISgvooBbhONg6Io5xgw2pWiK4I8TMHPdX73/1nYIoUVpbGdDGLPRLI1B
M6ciRa3eXYUf1Mic4Xf3213+G2WbC+kkiH4gg6IESobqZ/7qdJDHsKwHRgRMWLjT
chXQ595Wrskriy+z5/SwbfaTeMnfx5P/PfL7O1i7aOjFXnq5c3jUOAPts8LG561p
VXpSSSmQYE4xPgUoLmzlXE2tW1peMCz06HUkbHItXHYyT9jI/UdseEPRAjVQpDI/
bDYlOF+e53IorR9OJydU6BkY9qWIcnsEU4lBR9IIgdTSQW+BbZPpyzsPyCCs1tdA
CE78L9nCYceRWkppA6JJz4U9GQQoH6dw/TVx09dVw9F/tRCSuZARs6T1hCQftnnD
2rn7/nsr4UToXcQDCHFZPiLvr8NbcUyjUej/fzns1D+7k1vqLUUF7DcXgGMmUSe8
srCiPg4qath9Nx9Hfy/1uoL8CG5B3L6/Xc0QXjascKUO4rFZJ1dA54rNWtZB+NVo
ESC2piovOcucAJNBDvhGTY+0jhzh5pNVFPmHF8c4j+cBH8tbJRzDPD+XUtKLX+CD
UsexAVywjr1bQn4TNEWK29tBjzXnNMfgCBtBD4fEmIjEO877jGv9kAzcG+1EA9vM
6yx/O7g82vAv07dq/YY+sBpVDWrnqBZXZFq0qqrNbY4aWgl1v4Xw4l4+C0b1daAQ
0EXyVvSU9K3An/kNw6P7Gj8mF7/Bx2k8csjoDcNFeV4NsF1z/skpTHCWXxcdI2sK
mAG5gExVDCttUK5QDPt4LW2jN/KM24UOkY6Qd+FhmzijEGUv6BPxrOoWtISUS6a5
D2Ag7ukOKwN04VcdfCXI8gtp4wEdue7Fgik7nifrhSkSW2VCGEnyLRRiHD+VUYuG
RIDRnFPhl2LknfisISkRXX1gB+JcVoOTn0b87oMujZ/QUlVlSDH/oPU/oQLX/CUL
mEu858jFS1rUepicxHoXeTi3qa9QUgeVITj2H+JD2kEoPORP8l+JXG3+96jzSVol
Cks6vkPj+C0NDrgP4bVhZEi8xABusvW6RT7fNiXwAtOJVTg9hmsltaZPIhXyhZSx
oX3m9/J4fI71SHx+2QRSutaYgSErLnCfEeiwYYgbgNsEoq4xdn23QITm8E6coSb+
T35KiHNKDeHwL3czEtAh9WFTpm85vPfWZzWIfgLarX3V7fGd679g8Kw56WGG3F1x
o0BRAJtDCDMWgvIxtvLnUBCJMKmR0bpJLzHiUc5JljnwcXSsCzp3ltPOOuCjAHzt
IWj7bAdnfROrIfhHMasHBbeY4A2fkHra9f94Z5CZDshBvPL7liXnuuxwkIFeeE0y
y8gOxPwGee6g9umdmA9kA2f2KxaGi1HM5rcElJ3/Koz2MV7cZU+2qmRH668HPwDv
wp3iwlQyqnncyEAC/dVgL3IEeafbwEOgVBxB6txuxxKca1eSPaySpUBCN2j2z5KV
bpBRAzSJakA+bHk9ijIxjyXceh0gfpNuusYfUiZPIInVcMgJWonWINNsryKBj7pv
pq5ZBWEdnrrwk0K9qVZcNWdNWdkPPOzypqbCiciD4fVIvC4jeCkXf/QXT0qrsQ4V
08KEcOT8gVU6dSPFA42kIQaafopOGgRUiUh3JXOXoCiH4uF4rU7j6jHsNgSC5s4r
oj+9Q+b5UEHS7a/6RL5vFIVv8oAwtbrn6Py/nWkPflE+Ic2JOvSCjx529qyN2FHW
1w0tirgGJz8HVmrvm2fZN8t3pHL1BzkJn4mYGB54ATbW1NOlCfzUy1MaIZRkuYGX
jtSPSC5Iy1qQZqqLrqQEwxt4ntMONAjQ1PEuJ+3u7DWwrm+MJ02J2Q7lnLDdYA8c
Aosa0qn41LnLpOrvhtGr0Qft7rzpVCfSw1HbADfbR8JHAPPISvjn+yvyiOw8UGb4
YVdZ2FZ1PR77YUsMKJDFgvY3XXcqVxQWyM9l9EQP0AVyhG8gC5yGe0I50HIo8MAO
7cGgMHgN8vp//NMendmvCUQgYIJjm+aOulhK0j0oeEZcTw++YHRRlxQoK3O4CXQE
dD7XJwMVPDwGhfi3sRQD07AJlY3sEjysHMkGi9JyEon7y/GRJqKrBVBtUyqAfcF8
ffu46QX9sW1BINb1vneozWIH7Z5HKxC8q1vPbdm0wLBwOH1+7swB/OIYBQVznRkD
eIIzRxwPzUmoQIIVVQkkg6mcrNpNGeuZf01Avp5+wDgEXw+wPaMoK/4R32MLRrHz
4gzHGGAgCW6oIZ4i/WbFP07uDPzh9TqMYjp8LgusG+GIkeUiGV3ZRRihbSRoOs0W
BzHotkmDh3zBu2v6oNdq7XWdVzNc6jtP5N4GiMawagSZCAEdLc1wFd7IrPumZWdX
jHXPkHrb9LYOyxI4G57D2kq+jbcZMmtwrcRcefCFXNMZRmKgS9iwPml18X1HhyE2
j5bu3VMhRVcNMCjA74PUs03iyHh7YF/7szmymhFPQIYHl7sCUSIVnKpQr+TLU3RY
pEq6MNlu3LoiFIqkDP0J4jLgxFjq2kLdUQznOksfFyrIkCiDId4Me8Oct/W0lN+B
Y44Qd5xmW+sKZkVYb/8j41PmDL7CWYcHsZVNZszhKj78iblqEjMpagnOuNnfx/si
LWm/oU/ifH5W3C4m7sMY3PyQ74qP55ssoMdhg97h0UZgJFgBaA67bidNzXPnLEqc
EOAZEQv9I9JPf9bLq9qFra9Ky+ukdxb7grAMIhy866I2lCb6LX1zUjtTm7oWA6YR
T2heQMHLJObTSLUVvoSyoxJ0N9jNAvEs6ArAJd8IrjOdvbpSNfQFyfYyq0xXFfBM
d34VetE1Tih+FdE+MD+lFU3tx0Xsc7rIqSRt4zhKuy5hlYmJkk67RnfKcmACaVB5
qC/XgCYN5f3OhaqI63lzzsCXOHpDDQ6DviOICeXkAIz4SHW1+4qCPBrg+JL0N3Vn
sgMsyEp2pgruZC01aE7JGs4ny3ZgNIYqPqo3AHxCxkaZORLz/i1RoxuzI2XuGgdJ
bdCV0BQqSeMbpTVO3DEDd8pkNOF4ABMpZpbKu76epeBcd4ReC7oN0p97QMALH12M
rcY4ZIriYxhbJG2FCNBvud1r5+8sOVRUbPM2wc4hRdZYzS7d24+yJq6NfFuEJGrZ
lvAId7rMGsESO5zi6a6de1/kNtMajQ0q5cFGBK2Un/2N+5HlgCgtYgHVXq4YMvIH
2OQPKBcuulQOXy7CdjJNZpK4vGOGQUkj0YUzd1oNXIvf6i8TuIbGkNy+Ensr+tv/
z5GVPempHiWQHuA9BI6ACJtY9BPf/TyQubVWGdHGRL8du7jIi1e+LqQh4onVmjb4
dcdi0O0xkSyn6P3OvVSysMbyH4TsNXNqk/GXyHXofRJKQzWla+qxKBXOGIOHQhAd
4hq9QTdqnN0dfxMEkc73PABEA4n8uaDBVH+afIOFKpKE4kEndLkKzgZWz1Dm4eLZ
ASEUoJGslUj0mDtU0kF8Cp2rHVXaF13tl76KAocIGpeVlXdU2nU3+KUZM/j0Yw66
GhB4zfvi/AKVSpBVdo2z8XYiI46tyUvNucqSP/jQutC4BzZioOMyiw+cP9FDDzH8
s25vU0sqczPEYCgSNCG8USIwKXbl+LsllS/BvqPhOiKT8gW8Rqp6wp2M56hNAbRO
0BMmu97+Xz+twbWlnUf2YjYES/BANgzRo2C6lYeA9Fzxu3HzqHujd+QSZ+bbR1U4
X5ICCZogXSSVnyW5i0XdjBx2jOOd4fbBpcUbGKaPlk3URIuyfjwMk+arlqW81rag
LkT9DwgPjXIJTORYlOW3zDQYgCeVHbojfZBLiZ9PCHZbcls2+1HWblRVaQqvEFfh
F2S7Lx9fQAe9+dP94yrw/3BSZwKa/iEzQPiFFL2T/q4ViePqvCYiSBC3gLuV+Prx
xsNhJEJNiG0CLLe4JGh1trBn3MsatNLFy7MYC5WnV3UhVD5k7odw2iv8aXvwbAqI
7pxeiDo6BiywAav6Wgzu1KgPHE92tdZkJvDZZFxJSAFE6x31ANUIVy6bSppBC8yl
/wHOv+qx1Rr0DpNVBRhcB7ZdptRqiehgJGnKSS19V4wVgQb2GLOSQIEhwOzyv7qV
1dJ2ocpLJJ94vLFmb31B/EWk8730cjJJ0km0LlBUfXTVxT1otCFtD+p2LyH973ut
qXPDTchXNzlO5uUxZrntrttLhlPhCSL5I4lBsZ5j/Zgnim5RytJsnjoMKCqjmOUx
Z3r+ULJH/wjCKfcZDED1YAikSwZUxtWNmX1co20yjvc0v+esoazIfoCtsoQRDs7G
k8bJJV2JZeJarB/jjuW/BWuhc70vgzrYP68WA7FR63KUsTc8Qdfkokr2djDI54G4
j2oIXqJfWeGzbTQMn981730OkkEo03oW6u5UXx9GUqwFwfe/JKYCyqMqZu4eQo/i
fnCzejY2Ixp9Dv+Mv8oHHtUoDmJdJ3iieNgazkiSC0Oa13azYlC0lEUQCvaCeGIO
FcPM4QD+wbhcKdxF+uStgPKBYcXpHg4gkkZbdqDu7HoMC2PJzvIWFcqI1yfYPy7W
wsRCj582GYkKXL9WUOiViUaxvnQRhAlC9qMYmEsPst4s1Pu+xnKOmHD/5OI604Cy
U2Rn9jFvvsLmQ4VDjYr1YdUM/celBIgGa8qpPPXUZkuT3xWpy0uWKnYUzcFLTu0K
EfP2ECRw9jkYiT+LmvAQSxyW2g8jIdLyvty1DupPJONgdvLCP2riicTPtyMwzhN2
0Iia2MZuXQEn5O5aVxS264zb/w5UtVxA2zp2pirk86NFjZnsWzUSnMcyQSwGJxa2
Cw25PlKZmMsxPTZL8+va01Xu8iifkcWlcimh0bHiL0ECJbbw96z7wFKlwT7VH0Og
T4KFwsc2y1dabRoOrFudJVkcxHfRjcUfNz/rujGwZTrlZIMtXC0DErr46QpLKk1C
AibL6Gedez6aMYMfRw1BvDeR5NDakCpRKSa1zWkewvVtk1nfuGin0puSJVLP/JYB
gepJzyx3w/F0zkC7Rsgfuo4MxybX0l0kSYw21h75ecLz4xhD2Mn7Nowid9ZiG3Yq
8pOrzgDPT4E+zFUyN3NqK3X2U4QYImO1pMzvVQtnDVHrZ3P0bPQyo8hKLjgcAl5c
489Fp4Jnvb3GJANzoHYDYn3BVvSLfu2EPbQe5NZE5ragKwdnxU7BXRnHMWCP8RjD
j8zKa+eJLpx5kfS2j6qqLv6N9EyzLkAJqo6D2zAJH/yVDKAnRMYiuP4Rjogh0jsR
MTZWlScv85RhxLFeVbcfeDcfzc5+nBmy0jVPKoMSKXUrThiETraE0kkSFr7PwQrr
ZGCOdKTcjrOmivIT6IC0YTuFxD3VqPsj14crOJsi2iI/cQOdH6jMGdnAQHnCrp4R
X+J5SE8UGWDwyrjSnPRqjXTGO3cJjM8wqMKAlrE5Uk7zRl2FjCEYqJzD2jVNCRsP
+lb89+UunIItVuZntmCeuo6AwhZQvP/glq83AnCHZedpMp51wdaA4FERZ/GFMYg6
s3Z+9Ala2XG0z2MGkirvL1g+zmC5oC+fBbNu/Ljy9jWZqkypfxKlQb/0fOolpqL5
L0Z6kUyN4HFNxD5mXTeDiPwnGE1xQAI09t7nRaU5H8gUY3MS+qdASVGLthnbNgWf
9Fo+ntwbSvX5xVaVVGlWmQUpFo5CSUcIkSJyZschzqigdFHaCw3zzJj9z1Ip6QCI
xyMN322KAtDu9NIJa3o1gikMG9NZw2PO59KzW5iftpTh/kQqLL5XBz7jZM3KfgOp
MYXN41Nx+94DkNeAJ3NRsc80SKMJeC7ghrxjM81DuIBkS07FjnKg3Bo4ooiFrY4W
7b+K0FjUwFOUSldSZrZbwrReOPecJ0kGyK5JiW7Q83H8t2hzx2mdh8DyPfID13Xy
rEclq6xIjsXyjK07uHA8eYvX7OdzuASW3vYRq8fW+Y6mWAUxMmFMVBBqSCtOUpcq
gMR+2/uYLDj7AejZvtla4aGsILfT228pyW6z0Dax8BpC3KNXOExQD7dVtCnd035t
a6T43gw1EIixKw46srGBJIjbLwiibk0iLERrHp5lJi9ss8+JBI7V+dHXhH/bX0Lg
2EfgvAGkn3c9TDQ+SF4Br2hLYSWpRA+6LASS9Q3MeMdNCUrOAx9bn30nWtr9GDYf
nRQvlwIWIuhARLr/X+1KkMtVsP370PQX0C8ataqWYUG/0xo9WpxxfpzTGkJJ9lzJ
Yt3nBqRAZmNWYDEOwdHR941kNdJaOpeGLLOsi9IiEgoiZtCgwuGqfv1SfYSi1nKj
Pu9Izfw62q+eTsZ2LEHtukfmonH8RUivO39oLxRJ0U4d6hwSFCAFQOAG9F30iwQ8
0igfzh304caIKKX5ysROW4+jeIRuaXPksBgPkJirdEUvsT/vhZ2n0vvutgrQ8rTX
cy9ZgxmM1iPraaobOzfuygcfd25PTTbLjcjtXb6OA0qKPAwXGDS5IxlQBgisv7/W
kPthRQgN5h/4QsJiOHFvm1VeI1kg0UPweqZau5P62q803yqD0MqyOyOGyNwAsBXh
8Y4a+507bKh0u+ngFOPbVyWhN706WMXyWx2RgpztT78gmZPIgO+mBfXwroV3XT9L
zgrspA0+uU3lIAvb+R0R/OHkKZKDvFg1g5wpFY2beehQDSpOfsb6mIkz7YlW5tuW
awsltEmDZoLqaFHY/pQ5G/bTmofo7X/oJ2qsyZHIQkLejv7mquW7FKy7rg0mh70k
f930WGjy7auqc490QEh4sQl5XDkWGyjgivE68Uv2nqtyCRvvehIJPguyqvxcX2j7
XH71gybt7tLP8zg941lF/QuCLCTfimuVXdIECnqtZur7myp9XSw/Li6Zs+rDLv7H
sm/qoyH2UeHulywGyG1XG4VexVlfwePFjECdPSrjjPBI54SWwSnJ53LUPWYJ7c/i
FD1CLDjDOdNp+TV0fCiijGQ/fFrOoBTeBJfurgBy6+9oMJJ4Qi9H+LeUNISc0O+z
2dzCkPnK7vEs5hTCFKY4W3krCEKxzM/BjRjLQq2Pze8Hl59cGlsWSqwl0UPjpzdL
Ul33KZUTeX+i5bXrCy6xxkRSl11eWQIiSr+OOHAQSV35xhPm/qm7whcPYjE+dSIJ
C/OLNqLHl6vAY5yxO5vsBYV3FFdhXiTNwg9p2UVXi4JPQ9MQdcw+1E/85+VGHxTC
83CoRs/ugVc4pCyA7bnSzSjBgwPk4Oy4a77uFDFLjVzx/R0k1/ACgm0q4Vi7QMDA
cZR/oxjiVkMAz0ntS+Z84/i0KKoo0wbMU8KhJUzYE8KBrdh1jfj5+p6GNJ1gwhEI
9lN533OEX+z/T8LqBJIDTQLn/vjbxNwcrZaOVFF5jEKMejglYBZRfBWJOxXABBKu
TPhfvRKPsHND9a22D1FPGXtbTDAFQu79+CbIOl3eAvlJU5b8M1gIdQVjKBhJqGYr
vn0JGUmid38dnnGYIXGEiWLYMQ+IKSlPfPNPOz546IFEqOrYvIfk/rvQNHzMafGk
lkylI+O5pymsHIHkKSWU8e2+FG5KcJVSh/N5l3/PvHrt1cnVV+GjOAcblxQoe9Lv
OggVBj+WrEUM6g1CAopkg5Wurg+sxGctdlogKQlS6v97kMSLS/kYNeriniqqXOgB
rq0k8cm5tnyh1Q4HW2FaCvnm63qBuotL9hRe6MuM0C68/w+6uTGSikasimQUTMbc
oy+zk+dtT5SGNK8A+fBTd75Og0WK5015Lel++BRPykhzPJX1sKEStax2QxeKkw5f
y46XtMREcgzQPbEmfhbbpl92QJY2E+u/yybHTp8Hrj5l+CljnRQyxD2kG8TmIjYs
4AAoaqaqA3BicE7sjD76Dp9GQ/KQODKkPY7Qslb0OPRqOifQQsxQBmRIdlTlKT6B
E5t6BC2KngGYUP7ZIPGT/u8cYv0Nw+mOVAFmCDDe7T3f/6VADt1s71Z2NS6UMkYD
YRq8wKa/rKoeHq6c3xj9F2TjgSbmhpD9H5/6o9IFW1EcZgE3FS2RmA0BlOb+J/CK
jFImiAsLr2Yv7JXm3J5El/2rgvi4+0WWseZZZekgH/rR82cFEvtm723bGsrZhwKS
BHcFswzsnwZ4Swmv1bf/En03xYwr+f2q9XFNyWwbTcrUQzC571sHRi39Z5Q5BfAO
DrkFRo4mJvmgVqNC2FfI/EniplvFESVa5tng5oih6+a2bSR+wbs6hRfb3kaIEveA
8+0hVBEo9B7Ph5zOZTv7wis6QmWIO3nXGNRBg8jCLM0VVjo+BgcYCx2f2z2q7MBY
GnZfFVv721qGXEpB9vRGwcFIm5u7Rez43ZriSHPgRYrS26tb4t7DzSxBxYy+hDvN
9JY/sBJ5MEBp2He0mhEqgLz1Wr7GLb3LYBeSVkHA12LsqZ6KA1at8KvOg93WzSLf
4cDmOLBtWTeFZGnUQM8JOJL8cLkPErA+I+Dgjca7mnW45iLLv6rLcKczIFTUMaJZ
6cS99FnK5bPwY89zt4aapMHcYmQT8LHtlLENO79M1yxCj56EUs6e4mZYZEZyJoOR
CkclHEhub35zv+aGQA4C9HDOVAwvFPoW2d84CObCgitabyTE/E7ZmLGbD0gsh8SX
f0GlmvHnT3gZ5wILEB6hfISOLF637qQFzk6L388myMKhJLOYHt5YKpY6nBk9bf9l
WOr7mRDk9Pp4oJWmLRM3u0PUWILmiOWvuUxmbzD5HfOUmWtxjt3bkSEsT61fw0LX
uxfbWktll63MJ/vXj0pKmiWhjUwtOPZXW4WGpWqy4LY0SIEVBzTB5jctznlJz98b
rKGDiaqy2Zcr04kjihxh2guP0epsG/elhpEtS4zOYzx2YfcMLZC+YO3Fmr85dFOI
VYo90zAh5QA5y1ioJkKTTpP3Uw627ZrRsiIBgv9u4TaIcUrIH1AcW1Y3WCjk4Hul
qEyKfI+9iJZlhVMIkp8nVWb2UFzf3+o4nrYvI5wpGwtUSMKYEXqJNR8qaQoIgfNd
Vb7NkafPiR08T7QvP6fsUQqkVx32jWUEVgOXQwUP2iAIJVoROjDapYrlsUdue7FY
Ee+Yrj96z6IqfSu52iOrOJj+4KBUu5BLz0v6lvMfFGIx6AKeOHo0oP5b243NMW33
13mzFhqFwFAdXpIC1/0hDYilRaYs8UIplb7mxnPzq3YrofoOENcrgreEWUaNwYXp
/U83tahKDZm+2RGmvO5rusUlWQ3boXBipPkv26+Hc72kSBniakl5OJzH/pAXsVHJ
erfTzyvibFmvJfFADk7Wi6qnhc3swVZJbCx7Rt9rwvb+MnjRTl3qDP9Ng1r20ZPc
KAnBN//u2F7AgM9FMTYv+JhlAXnuCX/ZoOVuy04W6h3Rea2dYnooHSqXyNTtVGU9
GoYBBaF4oKdD9A+ziECHNxPdX5DHSOizWwAc2MVgfktS+zjxL/lY5xA7tJL9U9Pp
oknrUBvnJMlfXBCqqXldC6k1lwsOww8SR0sXCItdTe1PknDpVYQ7ONx1jal8shon
h3Wh4Ur7oPjGQv4tFYlgoW6dbbJDx4dvSH+suBASWBB9wH3ifpk6gqjBkRjPrBAz
8jp6jBp7cEPIOVWlTMBz1/itnIyX4mgDYW4JCDEpO2NL+4a3vUthQ0mZRxHDVxRJ
VgAg5fmC874lXQebPPJRLTQd5irjVPxQIvOMn83SO3ChNJZlfq+ehaz6e26kGaUZ
ry4huMbpssCbkRUHO5ivt938r4ypRX/t2DYliQJB1m3xKA+VxK+3TVUThvj/TUGb
CQqrABGF4QNLSVFjLxa3oyIFKx+NzQMZEBgtGPtXqfJ3TLJ5cJbLzH93GooStNOP
PYyN4Msrq4wdj/gJDJ1kK4DLlw//LMAaAoriKWd+8vIGO5n5Jic3pQVvcgCR+AsL
q0QzpWqi0GcTo/H6a+Y3arjnnUXf2/KFYP9zqm/2yxpz/0zRzpOE6hCXY8yXVOPR
n+lHwbSaN5jlATVvS/aPrTxbZybtikmiMi4r4DJj9K7XT+AGn51cg0m/hdU1hhAg
G4P9jVZfZvqqptOmQTVcu2c1aGLsMxSToAt4X+khZ38buMusgcj+k8AcdOfagPjd
LBoufR90wnkPU2LwE8nNeCb6gSJX21Dh+Yfimw53MYJ5QMZ2JBTcUhuhk3HLblWw
g0XSkd2GHC73ttTgwt1XQdbwsYNQkVxILt0qzaZ8nRAc/6tgYulNsexV1iSMBa7T
NvKSzf9nuXh86PH3yuTI1aN+yqWqLMG6Cw7Rd/5WtGBwk0xAMWJwez7V3UMmFwUP
KVMtcRQoqmFAtgzv9J0ADHcVfOCwPoy7L4UfstssbVWFMlSMVq/5f7u7rJRqtxEI
UoNGetoWAIQRvx/F3Ux1l110eNof0FJL5TRyeHqMpVSIUM706vBKvAUaI/HK8r3+
KPgA2geru4iXRKKRxuWo5G3HSaUz6+VeaDMfcG5YgUGkE6Hui7N1InhS5MUg6RoK
oFxMn7+2pSSFTWWVEngqUA0aztkrYmOC0Gj9e1iPu4Pyp2OKkqaihzr09Kqm8Ux/
QMJHkFofTuu6ecYvouJqlQvJFJaqhYt0lQJ5Oa/kGl0wwknv2UtIseT6kSh7ADOh
FQm2mYDjsfC9TSdm27ce57HJh9FSta7HsCWGeZprRC5APeN0L/fSPWszJGfAz97Q
SnxTBcIO6evpfV5IWQGQavvtrRv1xw1EWWEj0GClna45+A2NxI3aZGiH1i2Oe+sa
RK9o/vGhhKqyBlU5EBIK3wHTxNUZ+q1FjHZuzVllapkBQexfXqPl4x/5F9YU7ta0
I5NrQzf137ttpuTt2CDZITI97OVaYzQMFgVcYZxBrx0W+QJl7MqIIbelmy3lZfae
Th9quYgc+Ai8xLrv1uXpY6W8vuCR3b/d4E1Vvx4Sp41Cu5/X8nB5hPWomxcIaidF
WD/8oazZjPn6fVFtRbpLWzuef3LRVBVCH1zADAtKrS1aaxDtTN8fcVJ9ZL55r7i9
mAq2zX6GnTXbd2lq1r69WAdsvcqL4j0Z5Smxdz210zyotcQ2U+1vVOWEEB++6NCB
dV/aL3dzfsJhYq6VqPmBL20BMrNevD1y7IAf+VnyT5IHBaCndG9DVASp3rzsjbr/
R4gcZltW14YAx3N47vhxMo3YbjWNGfchw8bHx2US9ZMK5rQSNc7jBbLIhpmXcHgF
YMuEldWMWhpYZTS4RH1XryOpmLYN95GROfEWrVMfswbtJGb4pChyqOs7oOOAEpos
n4/O+ItnOTW9GFdPoAQhUYXyQHB7vfnUYjvbqKdylx2Ux1DE+gFWsQxHEfJ7EMuX
Sd74KhdsVR/AozEu1EW/7wEuU3oTQgrLUhzK+2d4kZS/wYpF4XkGvfT+nEkWDFmn
I8NMZE8VRcmA2sLIsJVtPyJeryu2KMyQN9HoO5sq9bqcXty3rjuNnL9tjg0xPaoa
AyoZhxe0eWW8keetkjEaHtrRLgVtCqBGL/l9bAUmMwWK3KeIb+t+xgS+PbSD5W0J
BOgBSP+D2wgDf18NSY4RHPO/ekceJ9I0VAndRlVk144LqsFM9QW5K6tczLFGjjgk
RfsAKzSZ3yWUzF6kdp7xxUw5ZP6AmemTrPRdS2btkMfZoc6bvujAtctwReC/hH2+
CpZLWiaaKWT4mIBA3oAzHRZzu4e0bxrXEY082hwdBXaiUmuEYUhfTXCNYK5wjcvx
iUwiC+lIqDEnWfcJCwFkhnEObkZX0I8+/El6+a39zFusXIb2y+5LKvUUZDAkjikd
K65tnG7rye/3DXn3VEpjgWlmB/dGUXstMJTqGMRqjeO30Zlr8pceDMqfQOMuUiXs
vAVnDY/NIkjFqVdwg/hwDyXV8AMT04Xjbtbzh2qLQhsNMgUcnkGhlxmAMf0bt8uR
fEE0XR1oEwaQOPF1o/NxsXDfPU5XwIq66Wm59RgInNO+AcroMLB+cNtUlInq/EZV
YM2I2S1MArHpg3nafxhW2HlTX8yfuK7LQiDD7mqrnL5XjRc6eOTmARpTR0MvH5up
ZInZmf9bRfGD0GeLi7/BoxqAs04Qu0hkfpHXFm1RCqu/h4O1DjTp0QY/Up8P1cTa
LdnnbwmkaZN3CcSu2/sMlxVTDVbdXuygqFQflQeMgvYK1fL75DkaWZ1q26gnkm6r
3lsbHpNTxwo1kM0aF6um6pouMUnkchWM9IX7CjBsWECdycxpwj6iwGoYYwyCIeXq
d9T04WidyNpvqLnQk3YBroIlU0uqOanRyF+f63DDnsB4j7Chtq2LtPH1F7gbMcBV
ZEHPTfZVZaEEkDCmXLGSlT/FruJnotjIL5tTy4IboX48PGaYcWy7PIKRqcXneEF+
RUdLjFv98xkQc6ywa9xX8CMtE9veqGNDjdY5Z4IgFcik6ZxIPfKU1sTWRCwGC61f
BvMFLjrJ5fD7NbFRDeD245WnGl0OFxMqnDUQf7EHLX9Oo4PmTRetdvIQPKCQWyzo
siknIdL6G0EwZbEHH5tRVbGK0FnYRmvo4D6iywqMApvWdLTioP7JeV6I1hW/EjwU
YsNwuy0XvGMNayyhOjrwGIcmN9Z8/M9XG11wvo+Lh0QCOfCFctaHhcdGk6mW5rVR
IekTvJ9B0HyECN44ZXQb5SkXSizqzKhA8ilSGSD+MiHhqfeTgnSm1J0UlZJRg/A8
FPZ0udhcPjchBuzMjPE68ObZURV4FdfewMdHyxT+YEyoigwiez8GM98NkPNJcYPA
72wgSu1AWn8kJOnH0wNYqNcyLADELbbnU2hzAAERt+LTVZAyGjOiLpVaAYpT4Ezg
e6DcqhCUl4wAJivuf2UCnvcFz7ZeeNaBDNIp6/e20ImrpJtxnT3o5uBZ+0wC2USq
UYxKMla5/bGeOPQ4L1ctgloWseWgPL9RH8YfnA18u61OZ5w5GYB1q5DgBf5K55Mf
vcEZmj3qq3OWj5Ic/xecsFzAIPjo1gUWpYNL2GCUwigy1oeGbf/WUbE0rAKaBwdz
EHEjADSQEAuOqpYWM49h1dlucfhJULFmE2JcrNZLKZQUc3z+h/g8eNHS2c/gJUjd
uStykwDo4THTtBw/yqL5PMa01g4C0r6zOt8s3ddvO/7xfskOqIzyaPWrfb3hMKcl
Gfk7TiGURaMavHF7g2/dnSaJdgEDcDeRhRtTkBKWVoVn4lltaj4/r/kS2tBBQhEd
Fm4XoQCUDqC7SGkFw5uKhvt3d+F2847dFejlMzekAk0wKyqJeTwJyVYgdVXicc3t
IRnXmU/4Hf1QGaYDdFWH2wkmUdAk6KgDzXgIUHHrinuXUqGW+NneSN3Vt2bl7Ksc
OnVZDFuPWSrJRDcYYEAGd0bMvHWVaQ+pWjP1ndI/g0gwrnaV+1rReojIDbdMi/qi
9zb1sxOqsNWsRA3CY2HijKlaGBRmGHWWFSSqgM8/3mpUF6npjEQivxg5lefXi8Oz
/1NTDuARs3re2agVR0Cf0QGj/NKNGWjYvzoynWbfm1czughAaLHP+TNd90xKw+bP
GpIWwjc46Otyjo5quNmR2uEZwFzKJt95X956MpGuWDHKUT3TOZ1qnQ+Vj1W3Mxdy
b4tO3OqUcQjfl4D4dg7RsL9KtuCpC77HUuDmTE4XzGO6W/FN9gRT38WrhnIMpZHD
mGxKpDUu9HvibEY/GTIMe65bggIupp17vvyDSAKJH3VuOTUheZ/jz2CHrl61WQ5o
ACH55IcSa+Bj0QAtuyqD+Qk3SyZdRmaW4P6T1OONM2taZXJs1ddzAgeMU+E+ZpuL
JwELC3/HRbfsLZmAVthWH0tdg1x5y1nH9Z5WswaJum8V4YvyFlCO7zQtSrVV02OO
KqxLlaCcAtCUD0+7xkGNfL3KJhIUc4we7XhLTwOC3SgNW4SntM1f1AFai/eC1ujq
IPtFrDBvbgV8KPfcIA8J8rJYGSVFLUX2OMitl6ubWu08lnUSYQi/1NgmtDwTtFg3
wQe6TXn1nrpkHjzCOksiBQpNv858YJCIKpXp0dRkvGOXe85aDsztWvKbaKAb9yie
ID7dZNM763tcHnb2IBs4CziggpcILQxu4Nt5xlR1Ick+8x3JgVPvq05inEka7CYW
iAk9bcomadNlGld8SHUglozS7xVgITzUyCrvZKET6sbQFlMOFxdpzDr/2kp6mBSh
AFeBlNKbFI0n8iSTj2pfOPuFCewr/VYykH+oHdI0Q5NIW3TVQQf1rAy3YZeWgvQZ
NGc38INtMXdUbMyU9GU8W0+hSjuVI9HRuDd+ZNwWEh2VaUztG6pKINv9k1/Z1SHV
ln5yhgA71cZSvzu9ezF89anFmHWj/eUJw4zjXF2wjMnos/NGc+nSWP8RE6zqms/x
esf4qpbOxKObfy+NRTHQOFomeRENcUdh8vZTJjuYC3knoeeWvxykSMyWG7Evuxhd
dJyi/JqKG30wloZvv1pw2Ms6Iy5oInJ9zTvfS3d/3pnQAE5SYqqBVk5RKSZvoKLI
hPN4gik8eRTHei/PwSDvPpSdqFD9gztCGi8rl6y3HksM2rjVGrLBowLebK9/y/W6
6NdSwQRh+d7xNPFmF7I6styf/n6pFqihhVwM2FmsPfTUp+W/RNztdssrwiidKvpC
jUPqqIChDnGzepAPlYhaWitoy9Ln5RHEQkEq0EXTI2areARW8CR8vOD4+6l8klI1
UjtITE08DQdAYkF6OFqN3FAySaxG4qs2/LXaPnQzlfmUmlDeUCFJ7LTjxjQXNdFW
9Oq9lUGenjIXPtEzMK+rJZnsvwQGeYfZ+36z1F/GRGjqj3mad90thuSMM/gNnAVD
cLidMP/nT9JKDCEfOBr2fPEo2dyk9hdPMv8JfMq8zacoFQuI9pwYuXMUtIaKOET4
akGa3W0IndH5VAKbAW3HL2GhV3tM+/dibcfZH9/JtbvmwIU64+Ab9wcEax6xC6k4
BCGXWOkq8Pxltv8AAOdMOzEhFqmiC+fOvEO0srzOrzI7gIOoA61D1Oo0+4o6ZE+K
CNQbe+HqjjM8EUxPzMO+FSOppLUEd3vMYKJ5DKC6/4agkGQV2WM4gL4Fk7iOMeVk
mgwfB6JBg00LvwWxiFzBgmsikEmj6XX84c7V9ZS3DtgoQrI33kqMO6eReWl0pQWv
KuvnwcCJqMge0PyI57HamlPEyhhbp1WEvE1+qfmvaVfZdhn7nJPNsAZVHLU6/IvC
FeLG40T9NCVZj1QlqGaMgKeOVqfsNehQ8Ta4ey5kLNwssTsrXBwMuphg9qUg6Sa6
fryxvhk26NX6dgZkuv120iq2nzXSnyIiqRMvpVcH13kVwbnQ47NEk/iW2pV7XD0l
ZOy+vNjRObBswQZ5eQkfUJ2XI46v9JMNkGbtUR7OEMy/9kaAmUhg+hXbW9TTjD8R
xyL1aiVqAz7EHuBqpS3os7x1y0Z3dsyFikcfFAn3ktjoChxFqaPikAK5k4DbN/0Y
F0ikWIeJkJBT1UolUj5avFrBj5aklEnB1Iy9a3y1SbXGTn/J+07atLebE3CNI+qH
BQi8yXZGzUwdomfYl2PCG/rRRqNXenDJtpJab+Ox+9zWcjRAmT1gWuGghr3vZmal
IOWvh9X2bQuniS32JZCgy7SzoU6/7+dDCHRdnPZ8AObgaDOwPPTh+bYylvFkcvKd
nRYtYOl9ROYNHYY/T3sfHeBBUBxh1QxtUpjWZ9HtsqwPr3SxaR7bPPz/cDk+roGi
Hp107ZaoWXCk8TbDCA5i57BiR1XaVTnAdXrzCt234/yk2W6CbTciEXqIStlhZZui
fsxvz+AxnDo3jMgUgGvgWt/7mS6X69FcU5dcakHmBWHS/5jil6npXvi/+hnUsslo
KiDOrj3KFPM4WtTf2A/GKmtCsCErQSS6y1lD40hMZVFmyDs/i1xUlNYyNYIPD4j4
LXz70oUVzkJ37N97mwxmzlFfKjwWcUgJtISI/5Ga1XuTdb51rd/NubM4TuUe3I4c
Oy+E2311J0iAzq2Vwr9SK//fr4UVh2k03+d/uoLesEqquyFaP1XWzzjWHKBc8OXK
ftoU4KPt1nyCCCswF7Afh9n0W44/l+Zc/lZWtRCNp4yVEjrjLAsAX6ZlM5BQRl1p
ci0Mb9SojVmf5eEoNYuEXrWf9zX1ONt9DVHYideDOD5h7OPU8t038h6H9zzfqvvp
+gsMLMZhiG/z5/73f6biFV4kyfSrIPZO6AjaulP+w0PnhEim3K0PeWrvTz+jW+vJ
uoQ8cm8PNT5Um9SoCH61gcM/rjWtH7M9AhEzTj7KY5v5Yq2e7T7FoFKk1P4Nr4FU
yOWybu7gtGP7wZgo3E/kev9lGRjxYvvoY85t3yyZTJKwMp85NBpnvclgtkSpE5MH
lnXhdEnstsA/wq/O4lK0OlbWi3CcAsChXg2UgJsLk1/uRnqHSzcbv4qD3lqnvTj1
YkEhCFEMGai0BO49uCkpUUGPYmnB+yyvxk3ZNtRV1JxYw4ITN63prDPpla59349p
hfJDIDgU0ETFm1inyJPWw65M/gVcyhFwfwzfcBTlaeohjZZm12CAXzjJMiAdl6ns
B/CkUtEpOGECknQqkw2OYxoeS+k4TVQQU/s4g6M4NlDa1HDy3trosLHhVGfRY7vh
FE+0RqCLlBkpnRYuEYubsjYwmn+r7Sd1JX0BqoeciWmeGp0OmA0EhYfrtX125gzh
gfBXFpIbiYcNBpcJypricEDuAD9SHO7wsCVg3TCZ4XKN0GpSG7O3ecOhhZOuLKLN
OrAS0UJv3R1OOMi1ouy1p9RsHmKq/7Noq80bvGloFVAsEqRUtz61bWWQ9D32387c
4pTBMPn3NofRjLCoe40skao6+J9GhUP6b6FsJRWnNY1ZS19DMeOGIAnbPWb0NjA1
Ljby0JUC4XXiyytkAXmGJbMWAeWgcimoQx602iNg6CdVPn0ClHwXK6w9KrvBIN9L
IRJo120Kvz7CpzzBDG8yOHLA2VpgbEumJ3G84a9XXTOPJeEc1ED5tThdqfTcucuK
Fm3XRyboJIS/eCw+CM3lMsTlAcC0kUhl3EfUYwt4AUQTq+TiLzFKHwcJ0EdzErmB
boW00Cvr9eLGeOPtaIH0S1Y5geXVpQdcnuywqUW/FV8tikQqLwPLmZmZbiJEppXV
PFjfw+C07IMdkxDySXPFd0eayKsxb0pL/4EAMdJaVV8fCWaWZ6U+d/34gOr+UilJ
vEiH5UHjNDp+r4CqycYfC/vk0B4b0xmC0daX/v9A2tYSxO1Asq86g+LutweNEWU9
sPEKfbCPZ6gu34xdqwZqIYNS0vbln7sE3oX3JZyCJcB01GEeXiVbe9ArvU3qMMFO
o3MXeWpHqTwLyD8we4LbfuZdHad/Y7RHbRH9fOK59CTUkIneHxKFCiINSZfoYeGr
qiUaYP7UHYKEPJeOPDXhHYjfDX0EvobWN4RoxnMcnt94gkoSbqhsBFvKF8PBvSwU
p0yazqdRuz35rasIXHkjCk8BQ/52my5Yt/VeYc6rVR7wLtSjz9s9uGUA1mEaZnt9
eCH8pynTGAtO5/ewHuQkotbdqaiyREgL9FUGEpWut2K/6gtJ7y08cx74pL3F3kf6
jw5JA4PXsKOiE9AirGEkYPP/aHTxGl5muz+uQUL0eQCfZhamSEp6opqB7M75naL1
Mmz51ed6hB55fzdr3mhf4tjgjGt1LzAoMSsXn/Fpg1jU3usmukj9ke7FHYTW8mO2
XTLaA8qL9bra91F+AUPfEuiohOwy/lklS8PQKgaHADbHoVK48GJMVAjsE3oZ4lPW
ykwow1z+6dab+WwiS/H3+sUg3VHOY9OjkkUw6I6yPModj+s+eVZmdmQ9pu/U+pKV
vfVvOcFoH12LwZzjGYrdxL4V1zfG1fDWzCJmpHQYewRL2u2XZ6Zde+lcgekJsf9A
m1FoYz8CfFMSmoLGYLOKdzdJ5GuOhb/OBPw8fN9M7OyO5tWMuZx6PleQV+SmwVBf
nFhmQjDbAUPHCv0hZG0yL6Db0QaMF4kT2zAQPr9yaOECBWWYIvk2YpibRRBjrPUw
9npDWOLZ1dVy2A1zFLCUzHcnE8CJaO1wOTT5d9jMElseK7sjgFLRY5Pk13VNWp3W
MCRNVD2TB1NKdoS2CQi8ruRAcSBPF2wjX5Btk71z4fvuaZj+ubDPWrHKniEyVZOu
GkpSoFVG9wk/KPsmgKxVaAphM4wjzFNk+HfJKC4ENtoK8N4vc4+cSkl3MdiCnRtP
pjuUdxLDVi+/tg2VDK4GPzGPW8F7Jb7GfZqYy6y6hlvkeB/Auaa/HQXrdneYbL7h
hXX69j+zexgboCghvO93MoCvh6o70oIG/UoX0Hi/IzpoaOAUapjiYjAceK7r8gao
ePvQimS0iMKkuJSCnoR8zLS8okbZcRHhPI/ClrinDHCCUtRGffAhAIM3SekRUmc0
U2hZplbN5HC+0doIgD5n711zPHZhXarSdtegszwC8Vu08k8alM/EfU+3F4RrPNAz
Iie2mlHnNTKit0oMtM5UZ+ZSFhALNRoLDGWAiXVr4hbW7CPoxi1QSi5KgctX7Z2V
qYKnlxxxULZ7nagAT5b0To1QEDf59XFV+GguT4PROXiptKSqVl2FCLFXjOSCguVX
IplS1cnBdaImXlgXBOI+6ICY4PMni/ATqJvVAN6eeqvMcFFUlQUgEDkUAUxbgbhy
5In5Jvt3w4IbpexgikPg95XTSDYCCXY/HWcSo1PoxzGZCyrTfPUu7ZLC8LWcPcZI
GQmAaQVNnDVpZi28kVBcNQ+k6Vm5jam84pCQohKDaraZHsDiskyvJY0nxfuLtxgb
s9ds5IvovUuFvizChA9ipM4Xi7JKV9RiLnMrY0mz8S5MejR0/VP79NK/EjHkiMlu
UiUxoR2xXappZ3qTHqdKrPdLCr1pWsNUvX9zIJW77/3S8bn8dR47RICC1wnULfHk
yWlQvFq0O2e8CizGBuVTg0TnpSVCCUmAlQUnybVilsNq7MWagvr/AIt2IzT+iPvy
o2wrQuBuDRdBJ3FaFLwKeYYku9o7neWPbxZa3G+viE+zoap79oZzDY5nglNAxoK1
LSw7YXTYMdbt7jVKlc3IZVd/DXNZ4DMhrOIxxA9XKr/IniwXhCHZzYhfjauv2Hoh
8tuBpMzgah9fdNiQzPHWqlVf9F/Mc/0+xkiSOJzlIUFB/AAROeimGhQMCwymBpcz
hbiZYL8W3tOtTN0Z+eIts+t2m4elqdAf7LkAY3lW403Zj6+RFBiiUPFP5Z7riDpc
cFAFYRO1LbX1UyA6Da7EXiKnCmMbZaqzVhNhVagdVhilGySrv4jUNw1EuEjlLpn6
BpRZ/25JtUhLxOFnrkhEC6xh5bin7pnpKShyOOkF03lXvO9t/d5sv5UdHBPG6luS
tfp3GZ7P+2WaHABLNP3t6orzOpMvZh3aMvqGBKjxVWrXelAt9HqaP8875dEF0pYc
1PYtTa37Ez4xdNwUxaPuJgQr50moIUuO0LMDgHaz/l3Xf/6C2L4ZP1XkylKsykq9
kq4SbDchpda0AUkunRDhJCHXbpNXZ5BGLtKOCBUTXHQCWbVHToGvkKB6uwLGaRx5
jkHltA+Z8mxq9F+moN6Jv/r87QjTMrwXfwR6H+9V3uAmg9NA4KcE66rdt96dufi6
ODKSAH1OEj+82vL1R8I4SwKqKZ37l25IShj3anHVGceW3BaXP0dAgmU8oKvjFmiC
QVMS4f3ZGVGDayYglNAQwjSzcVAFUWVhx3sSDBCYQuVVLjxb/44NdEUhhEMxYfU1
FRCw3aWV1urwTs0SOLFm+nk2WdggFv2AyeMNrVyq/JatOn6bMeqYXfGj6lyiHyFC
fWwK4m7Lt6EKMA8SSIJsUtWzG/UwpaU5UY9ugf75XbBuWEDL7aPKGR61JqapWQ01
3aCiiKpfnPNdH3DyffS6i0cxV98wxzCyjJSn6QZ/rajI0MOOjOBVENLsKzd5R/cf
SKUp7zUBfbhbUL2A5Bu7x8lDXfiGB3UWxsq21/j08seUwT74nfDx6z6606YVNtkD
m8J+JRitbCAt0/AJElaJUNnYwkxcpbgB1h9imdbTUO3wdayvZkzxyAnTDQcWtNlY
uN/8A2eX3GT9zGJZVLpPZtBOasgv4+HcSwVTrbJ4B7aXEuzIndorZg9fFiZ3aThT
NquJjuiC1ANE90d6ieDroNfsMpJLG4jsDqBxTqlWRZYAuxYVHj1JS81Z1IRnAPZT
6gSo5vP3xSadjMGZfUn00SPT63l/m062sivWHLQHtHeECWwMIoGWtxJbovDWV9Xy
ftUuRI6SRf+GzH/GM9nlIEMwq50ZyHjywO7T7KTmU/w1rXh9ZDeaQiZAoGe/J2ML
YES7aoRsN5woDR0m66UeoLbJLXGI22r7vrbtfuqeGmaQjRSbiitu+NEO5KH0FhzT
ZtbDbnhylfEmMJSFrURm9u3xsABNStqjiAKpdoX8PyHfQjXL5mgy3rnimU7xxlDo
I5NILMwdw6i5Ubpf2U8b7jxHT1woKPa1B7iDEzyxTmwZXvXwBRrzqW1w6xWfGnyf
AzYv/A8N+NoxrIJPwoUEdpEXZ5EcqqOYhk57qQwfqfKDrtvsGjQ2Pw58lvyg/Mpd
VbuiyplxeO0xbZCxUQT43SJT/oIxvcSQCnQevN1ZF8bMyDTll7u3w/88+dkXm17V
oXvhHQnM3mb7mq6W/n3Fza0ObZSedjbi/Pd7yjdUCpg95b9ywEPDmsWsspNugcz0
Je/qBTlvyeYC/XuFiMfo1NBRPgjrQ4obOROF449kOHNVZrX+mb7JDtr5RhHLbZ/L
4PoZcn9uvBk/FRMcfDlCcniUbEKRTHHcg5+c2BBKN2v/B1bFt1AdPIUtxD5dRkr8
op9UIqNECprp2Ogu3hLPlTnFzaLQFNbfwBuzxm3EiVDIRZCV+TYbryo/YZIBYxGT
sbPsI5SX+201ZZ31KC0Z/NDtFEoNXng2/JbxFyLxXYErpCEJAYkEPFp+wA0nxaEK
srrCa4OCeX4hwd6ybjirW2qUhgIHFnkB3CC+Ra4wHP8/SAf2fpTlo7xIfxEUOxqa
y/TpzKtzjbhx2Ibsmb3NvkkROUeWzVHfkbXcRQYVC5rwJRowX90yH1GtuhG3nVp7
9AK56bpAWsI8wibgaE6BBJsyaNYLoqYyaOJJR5GCmsX7MbPtor8CoAtOELmnlu6i
AvTmulRHQl5rrAkQHZ1fuGZIPQ6RGyEC4TcXw2pwapQrKyMbUWdNhbnhIFWF2cLc
7fRGNRftIYKTRNMWB0QBX6gDWP53UeRj3jhESw8nEs3GS7xJOFGkBJJVCMZL5ada
lujgHMyd2MFPaB3WNh2tisICocvXMv88vrehiICe32cGdX59xALLTH8AagQ8UUJf
6chNyJmxZuPw8tF3s71hGuezXylp+nYYw3ouq646ddxWkBzEmijpER/0KFF2Z33H
uiMjpEC4+up+7uhi9jPaX6ZiqZxZoJeya7hbqQQwGRbHBlwSPFDNsKUoD8+UxNWp
zXwtLG1Y5vPK/82zH7gWQgT0GH6BZ2fujI+pezp80AT0HJwC7Ps/L17il9LhC+nY
SpaBQHRkY0LI0zF+Ebbozs17dI/Hy052MTbiFwDmgk1MarOTHaJxaXkWKZex1yVM
QRgLk4Jxm/Lg2pe3IXjpx6pRhycDV9wPUh6mFW6S6UGnvZegDNe3MkLwzho/yxGO
1AmAT+S45KqSBdXD2ExCEjy1i/K6xcOPmSKs+Xzc+CADMr3I00VR1QWBNOUMbs/5
U9BtC+O6Gl+0yiUXFvVOcqOiZN/QiyVA50Um8hlnJFrN7BBNRAjY8NHH9cbhlAO7
gMFU52zZXgWyCE/c+2YF9T7P3F9XVdnh0B54+sMagOtgqfs+C4boT0c2PtQJV8Jv
dTSs1+h9sbalmXY/besgI+Ci8/LkngsK5YDwJp+4UUnHik9bqpqYnVsVGxtYoqBn
EJaIXHjmYTC/EMCTBUKShksIUkzWLlfqlg44GIAu58AMVlNTOvnz7gR1g2OIF5xM
AK2SN+Lqpz2PjHYo7rF8UthlBHRecLeaIlRACPJGXPhjiTasOCjrmldksFx6h8K4
Yk0PaZLaMl5PFAKxY/tKo+FxnhL9i2+TB+v4Cp54BdlgDTesNjYiVNqekJSs6PS6
xiC8cTqw26wbI9NcFdyCm8y0NaTcx1WLT8SfnELubqJvgjnIcRG6SAnyAxZnlnaT
tQn9AFRXtu06apePH+CgGCXLsk6dmNtF9H39spVgHauKQXwuIkiAGYzr3/2m4npd
j/jseYtg+C04BLULLXOXp6I6wYr5/6IZmqFC9Kv120ASJcKeYpnqpbLsV/iWqXci
NmCCyTclRzrH2FcsrbEgIh2KN0vwl8qypt/PUX4XsTocom1wrWlOz4A4lRKJ9rSa
9B2EoZJsI3zO+QfPOKa9CEmdlDTIVXycqgcC1T/TOR1zh975qcur2/s8aOsYq99H
MTZmCzya+JyOddQU1qbeVIjbX2tgFg8hmRU1tvm1J+PONocjuHrdiAF2mZ3lPSqH
kkf8xEpg+QY3+0cTLN20PJSqnJQz1aSfx3dvybQSfCpJgMgEVSajLzeH9yY/AmT5
8XnbkBSNkbAmex0BwxhLr5GviyEc6xf3VctBP7H/8Wzvt5zRjGDRzZqq9ou4D6DJ
UJf3RHBHTcI7L8wV5JRl9ezMSdfMQ6+glCzXB8LagNlJ8rqMI4hzSGzYAismcPPm
tpDgdZy6cjL/2Mhjz/J2r5hC9wtSg/XNNgfll/mEqDNjxsztvBQGwyjx5vFWwdIa
mzgVbdyX865vzF7jFqkvlVatwWn1zPiSm+81rq4jK2kRq45MZAMF6a4b5FYl+Yf7
PbylxCBYkxG4l3iWD8fkTUi+fBLaqovxG43DmzOTLazL7CILmZ8yR+Cc+VVgSmm9
2UiIdOgBYaLBnbCUvid9HVP37ogoxOfiW3PGD0LmrR7QeYbEKrKVRpaYLnfvcojC
pyArVf+1z/DH0TPYTvML1CDFy/EP0lmw42y9z6pTjLIIkgaWDy7wR9S9HCZHr17t
2paRmkLCnvhP9sMb5AANtlrI5rIqY+qewsH4HMqoFLEH04aaeVz8p9rzB3Aeh4vV
AKzq6MvmhZNezqPlkdCkH5v+B16MVPKha7UCOAvNFcbJbifrqv7kYMgyo9q50FXr
xoene0ICDnqyqY+VITsa3NGVGZ5vA7o20kIkkGkXQNAG9YYwgKD3gW6w56C6ie3Z
Mo3oS9XreBcnhFtkP+FRZhx8QH/qFD1i2Ra+/qpz2/+v+gicOip6G8QHzIvjtwVj
gvKSgqNeGvuvdyCshuGrtGplwglNh0F63uRp27h0EKclkCrXCfoTsi7/yesilGlP
nywERu/tQ9KrUxRiNU6gkNKUiS5r7e+jNpBqcbbpzt6PbM3SFDeJ026roiooB/63
kdJllRXYNf6vDRHBQcoMeFeeJdSTqD0GEByzlDvxNQygVQ/wCYDvzxUfEoFpArDx
2rju0JZZNNXpxxkNJ/w2Ra6sG2rFyvpk88VHqiB20w+yZsydOdjX5mOMpf0EuooO
HW5AaexHklRX9ep6JY7JHRLzl+a8uFFKR/oHT2wMLdMutHRkZFDUio138fGf+PHb
2DCaevxs302i/7BuJy+VP/3t70t0+ldMnoHW3HL9cINpagqXbnDIOsj5nP5yvA/H
TEzUl89VPYY+25SW3X7SChG1SjNgIAFJ2AYVX9dYdlNkAzgBlnfqMpPI5Tsx0LB2
+sE8JInNqTmotdgpgYCOiT/DQEwP5Ji8Y80KoJU7hjgrJ12DdBBK3qJT6tjRfZ44
Np/yqg3/oIutPw8cBYujOqrooKPt7z3wTjQc7Dop2FpZcM8d4TGZfZ1a8OEb+oBw
7P0XXB5LKwqhF5yBaEXCcV9IUq7hSEOA2vAdAVslN5eK6aPZajwnPyszN5Kzs1bs
/B53CtLS64Qq+6kPRLd7l5OmE/ICGUQPMOTk3lVlmlpaXO5TLBJ8YBd/08FZM1WU
bjiDxxmJj8AP0hyfHuEn3oFm5xMk4zI6B0tXrBZJP5g5zVOeXiil9N+pexEYqVur
UqtVOjmejuZvtZQ7/Kc6LbNjHOmJffP4wPduqQSqCUyeJhVPQviMURbgogL3TndQ
L3wWaHQwvkje9nlARsLBXXMJ3SrJPMXVCwtpY2h7tcJo9O10rF9y/s1cFjIzfqQf
oPrSZshKKRI2qCAtyTzxQ49glUtZ59BZ3WCWmNN5D7QTIRtnqLeOQsepMhpyjJbD
aN6K9agx4Pfj3piT0xriVEUmNHHTjNHRdWwHyvcL0OA7vws0n5wZF2s2qdWcM6Bt
fQFoCbUP9bnRZVUF5h0ec76Im6WxbD6Gpaw4YfzJthnGQayMGA8oqCElp6PTyWKW
FSsLrzP/ArFYK9rXX56QIZ7MkIHx035nK+XG2Lk6I5D1j3CbIdsWB8IAwY+6fPyV
1YlPUYuR3NLfUYEI/PXJG1Lvs/8/bvtdcTygX9zNiheb6mW8JVZdfw8ea4yjFKQz
1VuE1woCNsSfFSlb/q7jYk7+K4felmVTw8yF5Hlie0y29HdoL0E42D2j6JP7hNYn
4g3V2wYhzUOcPa1aojm95c04fNmQVgwxPofznn0VA4YwCJUXTeLmeHtT691pkgL8
uCmfhXfKV4/T1cqhFt6KezWHYt6CRj0KIrnpzdomCD0f79rFkU5GaVKPI31HIvQU
z9BSmjs9PTMbslba2o2QhWZ3WHJoc/vy3Lrn8ncTXId3iyrkZsuJXsJKRS0WE8E1
oHCrtHGDscEmj2RdMgzz2xS2KsIDDLJHojE8Je5eC/v6bDJxxS8NC/CJCih0YDtw
3MjjR2dOmMEmIx8RlA6v/rFeiAE+UVgXIE8LRwCpIvq7VqMv2VBH6P/AGuTR8TcT
/xrsk5LH5no8xybo/FlFr3CDxncx04k4gw/GXrvsaaBekUEjxwsNrzH0m6Ndhmc1
08t4aceRW7gNKj4+/AV4b9T5JsbbUODdDF8TvPiJ9rl7IKOASU1LUOvktcZdjXve
nHJGRdV2dT8JnAeAM93cKSgYDYq5pFldxC3+Puke6QGGGUNBSJqF49zf8gy4gOBt
gocE3fi3dAhFV7sfJyoAzy0wFJ8VoIthkVYn6QOXwCa+8rOJ73K597c49JqHoimA
+aD73n6Zr2MtuEIaC75U7TM9nTLHY4jvWFxw2Lb9JA4cxu3ydcYH8htwboh2qmnK
UEZYbGep4begts5jukNF5op2g0dlKrDqScxaQ++vlzolEnoSbgXiKesvbtr0cNXh
jqKNpQ7uZx8pnl665ZBexCrz6yta44ubCUyLsVMXG5VlxzfzG9PY7iFjzSFU2l8B
BHpSJxjOmsgOBMdhElk4g6s5Si4TI8xd2mlAFVBwEENHehJsFZFt3tgS80gwmA1k
yevrde0q1Y4C1K23p4Yu0haxM5H9LBEONkviZPY/OI4dzPID7hl9Kbxqknqnwbfa
dJ/1lTv7Y7+YlDs8pv0e8DhNR+vzWN8ktO68eZCK3qaVU0pUsR0vgkUFwSUyCYu/
WR7+m5vfcto0+zMUWeA162gu44fJVhVVvq6FQCqXcpi+QgN67N8EcO/jdPoX97cH
Ry/cwBPW5YUOpAW3W7mZ33mRhbENTI3GhUtRAjsHhp+IuswNMRDMM80SAjnSCDH+
qJaDs9EA/Cw8xxVYfFmK5dVQ5is+9+Yq5s7WqOXnNgMs9cMBzoSuRopvo0J6CmR5
8WrLIFhI5q2kfMjs7WX0Q7PEACYErJC9Zsei/WprE+3wM9UU+e2W1G4SPhg4VCOx
76eUsT+LDuzvwKyncOaBlOFCDNKic4Fkf5ocVaqWeWaQoM7dnSdiZ0wAePs1CfR/
Yu4yiY7UmjcrKzm+iLINKWkYy7HDLTEZG8iTtvsikQBEnepotYVoySACIlRksOhz
sbBOOiON/HYZ0JnLDruldEFu8KWKj70+P5hajXiuQW6NMtgFYFxwXFXATQXSzac2
6PiU8cqNtpsGavmKpQFvqcckG5C0yk4zv748A6qsQziTJkkiol/UXXUY/MUAMf5S
qXBfyMpvwKxtOH0oJ4lMitbZsB7STFrXEUteR3A3QVFSXm2mf9Gsr4SNuqVkwTQ/
O5LXfh/echTdSgwRpvIniNQki33pM0NgGjyuDyYi6xPHmG4AzPFlGGdDIu0cztk+
tZbRFIW7vxdD/B3cob/OWqnVAk62rmjNiQ8NfLeAn4DgUb/2MkpJM9ZQoIKw1xoQ
teinNAWV/eKzhybJyA7Arkfyt4nKeGb5FU9X93Kml+mj0+QnrloiFBJFw3oifcDl
tzN5oF5gRMlOBcHdYf5HCka38SRfoAnMAbt0I29vnfASu0XjqCcTeppEjYutFpqV
qELYud4neg0RXNeD3P9zZ+9ITCgYByjWsudQ0QD1O9PG/neMyhj8qb2jSSARng3B
kq1z8+AcsaaW3/BRialfVzMYnqle71AxnX/lcbAIklyJYGD75gD4x5GSaTDtJAyW
8oGDNnQFlC74/MrB+Qy62NwkXtYMm7Fl66ptJtAiule6YSdOKdbexY1tHvkgAqSQ
GlZVkieln8dXHqA8zPCRWThk2CwtF9W+P7a5CBp3DQXIHrPkvrpOzMdVwx3hCFqk
WoWTM07RBUpDjpe0m/DmQGj2QgX9Dtv0GkXTs7rYHo+HqiL+Jiw4LTPWuwMXhw6N
7L4Df23PE9N5iuHp0r8xrvsLhv8/v2f2gGAYg6SBPofafWcYaU6jQ/jXoGKyJNnU
DwStTSVWWeOSH2YUN4llaRYv74P3AWXQu0hpzd9u3hicr9vAUVzAs9gEmK1VBc8a
E+W2/v+kk7NiicRD5/WUi3Ka/EPjXpOm2Qrde/1Rbb56PvTTeTk+PH0rDl+twaVa
kqqCS4gUwTiqLKzDNKdwEeOud7N6idx96U0khFiaqT6ibxbrDMK9MySJkci8/Mvr
gebw+YbS2X4sUcXzTMZpOgALm+TalvlUUfbQnh7YpoMLqzYnIJQqO3IjF/7WyMgi
0pMQGs0MYimGKNL9w1CksvE+UfaOy9hUP5zjLSzOnBzJyGsKu19m6DW7gwb4lKJ5
2USkXN6IpQuYpRO7Me5Qc6gr8rUcFDNyvbF/0iHAeuDLsZ+Wt2Iil/FLXTuKM8yn
A8IpU1pwGjSpQXcZE2YF2HSq7isbaEQNfuL5vQW6hU5swkrek0Ekmy0iawhEC8H3
GVEgxUGsIBrRegZdsNGImdR2UlOOX4EjgNASX5tN5eZAkZE8ydOji4s8txoA872P
JcW/u0NoKt5JW5oHaQT3rrAEt/RnvSm/DQssvoTvnAZLBmjHk8f9aqqGfHZFlGpu
O77JDeFW5wrCW5IWTpplRwfFjgCBaN0Ywl6cXxWbHw89Ld+tue4IQWT40rcWI9+E
+hBllFAokt7Svz76/OIhozPxIA2qjR5ccYdlJS+M0axCoTCEli/ZmryjrGSDNzNS
6aTFEKAC9g5aP1E8hBfDAeKGXGjcKWVjo2bSfdmG6ZY3KMETHibh/bMEkmpK4N6X
1+I6wQt52z5g3vL3e7lr8REblMTfmPuwzkLaRP8fnNN9qLSZnUvS1GR3+QxGeoff
YHL88Cul1Bzf1TyuaMDkKK6D+kejK4dBbLvN4D7y6l+LAIiZhRYoaHRsJvj6rp7I
28y41fLV8b3Jezy/UAftiWKikVofrrS1p3ECdHEaPexAso6piMYF96QHHLTiZvJE
e9vnmGBmVGu3TQtJca2au6Zs9FHT6sI056VxHkAzi50vUpb2UwmLaSKdf5suaqvQ
4KfZ2t1s8vwSh8zcqeIiZwSakTFBo4Qdi366WmVM3iNXVLSBwm2c2fFxTjkIGh+j
7ONRWDMbFDW/eqy1Pg6FazwBOnA6GBIdzgDxR8aSWIjv2DB/Ju0G3xQNqOtl18gY
vGI6SsDA9JiHVKbqlEpAYLfLbt9kl6QCQo20Iuty08SZ7dzZEQn0QHXrL+qpmPpb
810TiY44Qff0zFakW32WKn6or+HH5kCvzc8RC/U37u2S0KcZyJsNW+OTU1Q/veth
fMvObuBTultTbhPDuEj0GaJayLsAbOizjKK8vhnPp/4pXt7TpxvDmUW7wpN8IE3x
7Wo9zgor1mVhFmIi8QF+7jz8trlKcnsoQ0bjD5P6O0w2b/6a1oAcctH9qnPWtXXB
oEyeqqlp8nrMax/3gJSFR4fnQaypWLXEuTwbAbG/N7C8UEcIBouVpj9sCJZH8xSY
MFUw8ke2SbMcpWsOHnd7bPm10PbtIRrmAam5sApJQZ/Z92rXMVRAPDIkbUVypXos
VNEJA2SefOVQor9WF1RiLDaBwqYNYyKisiSWief+MwBG7lq5OV0Kbue7t2sJO4X7
5CHviTWkhbIBe+CJqobUmPo+/6ecpiWiQ1KO9aT1vSJb/yt8pUP0fisnkt5YuoRN
K8O48h8mTs3nFBE8ua/3oQFiTPIlywHWDZ2HNZZCj1CbQzCVM9pFk4GO0Ug1dmI5
+YPwPXjwtS+ZJPdBQSOOexEdjri/rPRDhCOA6SQd8GIUcar95mK3sxXSA7oby/PS
yr+mxUQj3redRnqJ4COArOhXng6fAJffreFLg7HZErPVRyvtD1S9oAGzQCpTtTK0
dn0YadZN352oX1afBcIzgEaY+mkNH+VfmsKLMJZR6XZS+oWAqeR7o1NQWSHxTnlp
+huTlRordeBgoyrEw2Wj/M9MtJYWZucSeSO0CGlNCgoLXITOpX5m57phewEZ69zf
+F9C1/hqBuP9dHIbI3LN0a2MipYxKv9+YxIKWS9hIMSz5YCETIyViL0vh+JUh887
DrBCe3c+sWzncrVUa/kv2gJUAxs9JEJxhg1kI/ntLCYrOq/lvfZi2ebWPtlXg4bS
pBCb+UoQ1SWguQjfkQa8OziymHq16i3PAt0/2GpvewOv5w3MnOV2z/SzkleRAoPe
3AUr3xS8xMZFcMrX5MGJxnyL5d/10dEVRpm1skJN1tLc0nP0W80++KBFXjO6siGx
s27uMnRAEc5iTE+ISN1ZhvOFpzK3YqUMtlSuIkJ9Ufk69DyxGpZB/i2jEyl35vtT
dSjsnG1T4p9ESWqNRPZGQnbt2MzF9mvkWIyiqUlUVpZrbUvREZsgqW6cVVXYKJ6a
o0byFWKlrMvxV0kt6W19gd6CKqGV7fqAgI73YHLcvh1+XWZ7Neu41qu/RMWcIkNp
xsBkTezrL8a02wPLUrbZ7H/QUJUfju2jW2FLpviTyBNEXKvlyP/CKv3/XfbjoMPZ
w/n7CX5OzTsIuGUbyuBSytzwX5jrkxq18PxYvNi5xLXHeKeo3WqX6XHlKVSyTLJ2
UZVW2iuwu1e45stw2nDrIX2v6SMNS86C6+JUauq4TnIXIpq3dIJIWqqwZWTiqTtZ
srQT9NcWfvYxYx/bl2+NMYvp3y+TKrcuStxG/J3lJ76IMFfhwTKMySHyvJuQ7Z1k
/JzEII/Q1pxejb2YCxRoVRnUwbUZuMRyq2Caa7dWrWOjXwbzeYK6t8ZUoK4DWL2R
3XSAdXQFBGhm/7JOPp1SGI0AeiDgD0gi+fGyge1kbv50HZadiLW6jHMLZ7vBaLRf
Sf1kKq7LUuRaoMX7rEYJDR+WVMC2tOp5aRh5sgT0d/+wMNmWL1CY2t4j1ojiAUK+
2jvfGy1lsVFV5bTrnDDuYUTta4sZ3znAh2D9Uy+iZog1J2EZ1B+YFGMQgd5hichx
XQ4c3p+KedfZzjSyF9ctOGdjauegPZHLpyP0yMQ0OlHwgFBnwnX5LdW+uAZekBJx
jlveL3i4muVqne1xqOkoFWZMT6qEe1yKGR40u9nPyp2+oCsj8rf+OcbjlxGa8qrt
nYaBVK1kCQ0QCZVhToMV+7GG0G5eHyfBEnNrJ73fPbVlbaF5OYBt/m1f55cjCQo+
i8fVErBhgioc3BGMIi4+i4XY0W1Lx25G6O2wA9HFLF18JyEWitrCJicVJLqEr939
35PWhYGWn53TvOy8EBzcE8+777suYQ+BcawhdJYpzF0Qr3howGSMEgGN1k6oa3rB
2gZIaHZ3BtgG8bbScpD6+lfnijhGoVmTXn+Z599IrXq+hkgg2DAAdzRcsRkHSitg
czFc/uyhd0CNpNwYdqwnTd6tbz2d+UKMhVQchjnU9dFGNKjZ1ibiHt87qDsMigJw
aQwj18s0SrjTgpkJZU9A++bUCx0RyFgGCZn5cuN2O5s/RVnMBSh0Cv54q4lYMdj+
/fM9jRYPiIgseAdbCtUblzslElRHDZn8TFKxPGi8MrGgPv+2q4jjw8+dy/Htotz+
YDlroA/Lk6/WUSZMRIK92aZjZN0HK2VvkNazO6yU6OkX0jvG0UYWFZDVbLW1EEtz
WeS5f2AahSoyDulw2jqia+wwIUpMLclTofBSkFmsOnKZZvS2Kn3DzVDJpKaxOV5C
VyUxmHkQatqtkyC14a9KqYRzsi1eCOkj3e9wF07kjhNxxZJ6hOv3NDZyh5fBo6lc
Q8xfZXwDmug87RMgcIYJzUOl23pFyBVmwUEmnNrXR8rrO+mVg0dV1+UknQ1g76Vo
5Yn+attzFjqHJpjcH/hYrs57BoV4nhAwSbFpszzHJGyb6fTRxU80I81lPWCTL/Uj
8aJiLOd8pYJLMb+UZI6CtupWqLaot9cL4/txJpKfL4vhhIEc1aj1kaV/DbdQyf/g
RUtNDdKO2t7DDBwUWM5rhPEwmWS0wePB0S/TeCjQoVdxGCsk7S9J9IE5L/Lmrpyc
I+/mhih4jpNcBzVkFtHy9iAGKEEs4B5fPlpMzBN/0N1nFneEU6HgatQi1PVTVOak
AdC72EZoRw8wgWAC+SGeeD+y5xU9JHso6aBe03QhY9ffzaDBfbf5z4ISJK8rcliO
CtUmJOOZgapTXZTrQWd9txKlaHbAjXfKi57akFxqWnO/5hOFm0KVwO+u1HAFPqVw
+V/QXo+apqnM93h4XdCzszs0d36jmLPbfQE31JyIe+7BWctq3wvnDeqTKyzWzfs7
yOih2oh78gcd3fqxewTkqcJDbUWry+tULV9jWbPLzkt5lWOsUaAINYIlvDQoWFOy
nFSIIOSHjOak1saqsD1LVtplH13MiSK3NqM1WXsMcVojQpkn4f8eUZq1bc1+etQe
evaA5OpBSi9hsgvNGXK5j53epqruNrg9QWtYg5AY3Up8RNnycaoZyjJHyjAGz4cq
j4Zf6Cczd1G3+ffEG4Gyi9bZIiht4cm5OITie7/5nHCOU+c0VXOKwnxyiHy/bD3M
AfxNRzds1yWOj8yPStylbsa6NFSxlEcZDmO3mf9ACY8Jq7g9hHBYBF4w4PfhtfUZ
mIdFwSyHqy2qmOy99tAe4I3SF28cI7XMn0tKB70E5cwws16fr2xtKRmiNrEBJsHR
A4JmZeAkGzpo6Da1HxY439CfOeoxLi9y3iyD/eXawGDuw9JvZ9NllI1XmabGHm0e
bVmDeDnlmuTbTkObaPALLoFntQMFIkcoGD3272R1QjWKoWuJ4ybzIuekKw74wN/0
J/DBIxNI6W25H1v15sT+yGkiYbfw0FK7kkBigIyyY9ZvgXSOv7dq39TWKJMXn/nl
mCl3wTwPxnf+jMY9X1yfJ3nwB9rxUt8qV3QejXmZvDimVwkcCMQickK/oHlLsoxA
MY7U/YYe3yXVevvr082emFu6B79cmY/CEBjJFwlwPXXc9h4CnkWfynTf6SkC+ekn
vf25EalstAqoOO4K/YKR3H+7hAdBY5FDWeDSebqnBgR6sC7yrT8yotDl8QTt31eM
dGmqW5cvbyFyoACOLtfgBl6SLqMvhNwzEsJQ/vC6MWHYEgS5hlCYqhmzinT23wSc
TUuR4/YrL/jKkwk09AgkhNozOBoSQ1Jhu+TWLdCRJyvXBJrYn2p1l+K/oL9VkYP/
KFTsL+2FmP3BS1hjocApn6PaHwgoor3YHr1eYbTJ9aKD6Sdo3vPhWlxn3+UT9Ndf
4+Z8Ki63FRgIhC5FAimBNeAUkG+1tix2JOpvQfAcIGn8mgUo1VfMqzHHazFus7BN
L6QBe9w+9zfZdhifv39xC9jCG+nDTF6c9VPEaDrplbSbg4EFaO4IaZAld8aSCoYI
CYA3aVR14GDzEJ/U42Tjr1L0MXllnsx65sLBojASyrqtZyna9nmJyiWrLhgkqZnj
nKk+pcAGelyv2Df8tk9IoLKt9isQ9KD/5wkoqTz7AmFfu3+/3bl/ahZEX9FCga37
ncFH1q9TnlagGTk0EQEThS8TAW4S5dFduy76sf0cjdS7iwo/igBcRpZRq17zVTLI
/ug9IY/i8u7Y1n+09EkyQyznP+EH7T4ObpGYuEjKo3hIhQyq4zp/l7QNd1ioEnBQ
lRR3/JoVn+bb3asto5zyaEr/sp3zUIwXKgP62oqlvLiIfz6qtSc0vNzPhtzqNS5L
x/LrRe3XFuLBHsmKjIiCIhY4gfqh8DpPDuPO9zeGFsCp/AVNjh23bX53dOHG9427
tYs5GFwtt0BDxNyb0VoH9iyiaU+f5jHaLfFqcKEVJwupdzKDyXWrbgH+TUlLlVNV
fqxNUUKfQUkhXL2Wx6xaASckuetqjlkuZ2tH1L+SwGw+o9wvqRu+2bzJ207r+i2I
aZCo9A6myxdFiN/+KgUrQQY6TcGkFstGi7KvjYG6SkhIGAAdp3X6Ik2xop4OtnDF
uRGQ3SK+ndSCtvFQjHXpmuiJRJ6yLznUo7kiDaN0UZ/NMj7tw9cQPeqZaC4r29ch
t6nLJsGWnl26nMyuEmCdMZ4IMtp0wFzk0eLRPo1xXsWCu+2sizBvVuRDm59woffz
ACxVf8j7AzWc52py5G7IouKmLITHkHWCvtSdU6lxfxTQ8uGKZRHe+KlMD3c7M35R
lEgudamDnU6PyNitnNlzthuJF6zy6fCv+HO9MiGfHasXUJ6WJZKdorfQLORDVw00
ICZKvpbcscgFJ75ZNrz1zUtvPLBuA2W+nv+DQRQV+Yo7XCkiJWbXRJ49t3GbrrTF
Mc6UFTMXG8UuAUgN0BKwpl8suoSAdITcV72SgLH9CaTQC2KyYSr9E4AXHlqUJHOc
JLk0qTkC5BdIu+lQblW6tiBPSw3QHVZV3N/ec6edrsfZjZZyUyL1O7pX8o8y82BB
WGCB8R5QY26CaXVvKLkKke362uyl5EgrKRXjbRYaQ6sz952LzoOmdsFfPIkjwK1y
MJUbmgWZXzbDHticX+YEIIE/QZWIpvzBJR9jSzU6KCquQeKIfqNcczjO8HqncMMW
Y4e8kvnSGubzbnxF0+MDwR9J+9xFDPdQ9dLSQ1i5AX+LtU2LppkfYpf/K0/kdFtI
+0e67h2lJCh3RoUCzy17mS5geLWQIZzTvcwE3cXBkoaK7pXY18OIOAYl7Y4DwpdE
vqvmQ/VP7ISiPsZUJSQumlTKx5/10t0JqL7g2IDMFNN9BiVg4kW+4KBSYIycod+Z
cB33TyreuGvLWfhJpVFieBu4eMKWW6BdP5TXjsdWBRRCt9vBrH8sfhvuHcsr+vo4
lfuBCuYaNpyGp/Cdcw6Nck+8kUbRnuWUcn23+Lg7NXfKsGJ/UjH9BB4Btk+am86+
lQmiLwJ86Glf/crCj4nDGYneJyuugAIxN52ouEUEUzUZlCU3lvDn4xnQzqmKpr/S
SDymo3pygZa5POQETYlEhX/IAMuHVorZIMF2H9Onu9IImyTl85b+EP3EWl0brNfL
XJF719NQYaAX2D8XdF8pRxdTpc8xBDh9oEeF36pdWUg+Xi3k69aRYtjF5dOli72F
gevWrbIA7k7RG77FplMkKyPJEcKBtgGguEKddvOu27Mwz1NGLTsUxwtN9ws7tCNn
zUEpoc4Rlex3bWWsF5QbvwKideJ43SDCNJHqUrhX8Oj5Ci3yksHmFYy2esqCb5rg
Gs+MCbyhb36b/2/PaSa1lCJMA75W0o8MlPAqkdrXRpfL2P2/QRRYGJT7CGKFsGmO
xpjrbPazLdFK6Kdu98/qdNhiKtQYWGc9WPW3KCYNkm83kRm+lXgg6BW+MUWyb4ET
FSvCWc1H4lYZdNjD5+OML11256vi1oyPDYlWd6M1UHmbHcme2Y8kqpRF94WpQiZb
6Urb5fKBeZRhof4wxR9H1sKymrW5tNA6heLi0y6emx8UwlgxN8kAiDsf+K5DoKkC
RM3Dqrt76LLqnDfYqgJioL3iiBIuvosNSaDaY+TKnsp5IP1IRs+tAnuM4lLOavM6
90UgI1hM20Xh0mu15OAvm8X/I3MEwlYozZoPS+IdeNwbpxtJekllptd0OiFKWGNc
Bu7ROziND2u3ofdTB5g8hXtjO9ORgWOi61Rk3CbsOvDY+um+e4loBQf3OgcktzNU
KFxDMF175DGQjo2rfVNfPTOurQhQsjY/KG6DvSSwPlnzRlcTqxlyJbvCTL6BcYXk
Axge5Qcf1WMWmEiOVZf7d6vY4oQQbVDQj9KZNliM958/6VZBaGBfLasWcwJPneJJ
g4aW7mewMtad4WRtfJyQygO9zzlvy6eFFp6YAO+NX+P4HIzkHT7oHk+8vnUII3Aa
OVNasED53PN2pH9UIw7LaO23b3dP/yhrtj+j/KMQ6NK4beMP5bDV+g0kEv/7Oa9S
AlwmdJwbz2Foz4jDy4EdqM3HHBADaznkb07c0Cz2+wTNolhHlriDmmB5OAIbtMar
2w7gXxSYLpXrZTzySY4slm8TF6PwcStABNv62xihAevU3/hmwhBINMXmzBUxtXDm
rJnhvxTJUPbkai1C2ABbCNvt/PZJI1/xEZ4384Jr9caEAv0XSxU3eJKWDNYMHpU2
70ihTAKCu4+01u76zyJjbO/bjS1BAisE6SAaKkvDOiBemZffX2C1oZ70DmNEcgfg
zo5I6ZQVCcAHvXRu0MZnLUTm+PusD9tWNMzJqq/3MQLo5gjMpiNurLYu4c7MV8Hj
4lyh6I0bAaGTebu/vJfhbZCHNRXWw0GevoGofz4haq0wLZsjjVUJLrfHWcQkarpt
HHCd8n36yLlT4EgXyZOdHpbz+rdDQsAEhYw8AUtyw2bVPPVsX/wEWKnwjyX3DYUz
Fsb3zuQ8pq0ORWSx7jwotS9nDdw6hKV/FqC216magkV5J9bfB4LsSAjZCeqadRUt
Coa3ayY8j/oRmDCi7emwqYlB/F+9HR7rAVvo46t32ps4wpTfWJZ40Ub32EebQb99
5vOGF2conzaCnCZfYdsIX8CgAoBa7an1PQ2yg+NqvXvsIp4Fckki1/Rso5MNRANa
I3XXqPFVtX2n96Wwm6zt/Zh0lc9IrPRrro/MiJeWD8RKjVMqIQAN3+002ZmC1pha
lbDwoLsIlkgKWdu80KCy80QkA+L6ckH7QOruFq0QntaYgSZvEbGdpvNl0V5zsR26
Mwwz/6Vrwj9oQBISjL3nY7CR9lzb8RKaeJxBs2C/AKkSmIOryqrMiXziwP5+V2Y9
hhnMwuaSO+nmHbAwcQpB7ch+4c3bQVh1vVgt+7He4c7l2TGqRuLDqKl5wFmiyq3f
wW0hNAftrUPxcv1mRztP8Jxl5M0+pkZO1t/Jl5XAAgMZQZjEWRiwuGK5fKkvhlWU
pcc483n6RlLeDALocJd/p9QLP4YVw3WAMOvaf1bsgtnztnh1IMOwWi26Pkl3e6Jk
yO6fx2PqMmdLtkz8xZbYolLPW8WgZGBbKsttb80ntIcmt80OJK+RQYeQxw7UwUQC
g1gqgYE78TpTd5Ztb8PAIdMe/Ak2G0BMD9Bo6NteLCC4Icxpnn2Tcir7lhMuGfaX
hznh9oIuHg07/DYmxpTMSemcRxUbR2vSzwvXzwjcwAZFPmHgPPnyiOYqnMG0GJCm
zmdf8b7ArE/uf/pc0ZoDqRcO+dw7YaiVPSmaGuXHEmFylkn3c4XYdlrWhyQ/zB3r
URg7GgKmUn8rNhZJwnmE/Rf5KyRzJZlFTXwl93e4skEld5XwswyZLrs4CObOE4VD
GTmva3Z7feZvaOtwBxt7kSxGCb30J6ww+74P+5/+pyDxxEnQnneGSnxjvkk5RJfg
RMLJ/sTAYC7M69I+wYdASOzKBy/lUdWBosfP5/AHREkaL37+3lsirTyqf3pXHbGy
VzyThVwKhe2gz5NgfKPL7IJ6vMN1CGQtCUUnv0zFOMNaZ0Ci8RkNuy1kvXOngXgV
3+zO6yo4ad1iCpM56MLW+lQNTM/dYePGhbspM531LrV9429H8sWG+VI1copCyuMo
yjcZGDqHYJCCcU+u8BEbmEUfwfxAM3yYiZiV6TltEszSYX2z4yrNhw5cXiHk82mL
3accRVfys04pk1nJbxdEkIZ8HnMIkswW55vm5aVDC2VmEVKwrZtdz32dQjbNKfIE
3voCH2kPY04VuFjWc/qcur9D4wkcpUEYsDz6Mel9feXQF2fqUaOp/ou/QJSjC9D9
1lEdui46qK4vxF3cWCSTiQUQAzIZ4dE3HgNV5ejpsTugyisNtsyb47OU6nBTBgwc
Z8VhyVp4Z/gpcmu3DvgN9PEkvjn9Axm5sHVkXqSZ6+uHq3Zqwskrq4u2HDDamEkO
LUEZF+qHcjanLe/zKVTCQ0DYxwDoKvjFTOFlI+z6bUMuDgoC2LIROVUs1/HY7nBt
fJbnYu2mNtRX/431ca8W82vFGEgwTstnN7Ps33MbDwKRZr0EAP9pny3QsZaqRVDs
jv+JsAZ3HkOJIVtwhYgpQcrGlI4TtDFc7La0XPaIYWwMT0qSO6aiiJv/ktkmVq2n
/GvAYzLMxT0DxFanS6/LDIOfqbF3YAaw+Lcs6sDkzwC1BsIZsqlhLFZrmXd0GFPS
G3RQJa36rl4KQ4jfIdj1k3C/v8V2hPvSVhWtV4M5tdZvYkU3WDkhilSqQhRueKwy
x9BDg50vuK5fEhk2bDhRlKesIEm9ATM/TfUFJpdmRe8j+McaHQJMCor7RMWg6NOq
38yPV4f/stZRaAqEAvEByuYwYQHvuw+jhnWBvie5Emy2YLt5kIRi72NYuKY/l/gO
7VlikGym14sO64UCA3/Na4WuAewnQ4ruaItf2RYRyJ4piA4YU86T2MGTAin9YIQ1
ba3sabApe4bl2vd5rvNSC6kRLDXj4GPkHF9ra9dYxSAa1d9ycpSSjJDBsy4jHeCZ
tLuQo3fzZaxyowuNSIPuw3oMX/eSTg0/mEWroc3/7RvszGt2t4+o5oEU5f3G+ZlX
3zc43z5LOwjJE36GRy9tzGq3JCu8SiGEr9Akbe5mDTcPq7uyknSrS1Qc/zIsQLzc
e2w+FaL3gbWm/Ip+Wz4zn1HJPb9GB8nQxa8Pv8Zm6erFb4PmfANy3QVyoYBzW/Jy
/nq+efaCgIRjsUoMjsj9OgLNfP2j5IUhKanszMPlKAEwBAYMyD5bIv+T9Vec/8j8
D5FJqpkyHPm3RtLYL8KHgmh3xNeDwtE2671ahioryriSLizBiB6BPPGv3mbTgBmf
TFpLSEuC9hXVZ2zrNz0Fkg8FXylkeCQjLe2w/+vZU5w+NYrxi6OILwtNmtRvcq/i
6dlGn452DwlNyilFuyh8zDD+xpbr4YiqdnR5h6chxdXeNuI0Y6zlcKNsN4ALnC2L
4Eqa5vk3TjR8P/QlYIhQPtd+xduCh+OR0HQhm5i0G2cYFQKa0KZaLCB7iPzy0+9U
TcdkwRL0yYaOeJ7IrGfMfD83Qu8dawIGHJkHUpZhjsKMuyscwlTN5Tfp15Xj2RC1
4/742TfZTil6dkL634NMbWyxFnfdLnJ9EVL9NmSbVtJhOFE5pxB2sPJJ8hJlO1Bz
+ViCJE76tCplRXXjrR97TrNooDfRRkL17YRVqJSnOeIYe+RACVNKBolIE/PDcbdT
VJ4v2c0jDNn1wOuvcJUttb1fEA8PFiwA5Y3nSgo0x+5DJm3ZPBwGmWwkmpIgTyaQ
+O4q78XoweuYTbrwTSRrrV3q2ZM44GLSzt/rNTisAXRyaAvnnSXFUmXa8Ihl54qt
r7/27rJ5kCyujKQggdi5vtHPyYi3O/wrBheXINCljUsCES3mbWrUxKcOf6Z7hfJW
JwxAHeus9SlIttJoycTUgqebFv7MBi0UAaD6kIJ6mAumxMYTMM8WyA1jtqiOlcoW
T39ajkJRzMhdlf1vy897laTncFS0N6MxYEvxyVx7qQOhUMeJ0IXuwvj1ZgkC4ldK
x0To11JHWgww9xQwQegPvKDUwVG34NlLd1Y1VF02Wi4yr7Yp1yaLCXsjTLEp/G3H
J4y4U/v9ZTMjN4H0h6AmI4MlZeyY51WJi9q1Y0+cWq/oKaMd+821xNz6iC0rNwX2
bwNd1L8bPdVGOPgujmyNQa2gN+UB8Ik0prw4f2MtIGO9Kso+6zyJLDU0wXxMDGyb
RcSxjPuD9jsw4Ik53JlefPwhBQ4lMkGMhfKiGDV5iA8w0WJnoU37S532pX1U9g+a
iJ2tdE5sAtFELsNEZlWep7R61gqFLVBVv8pBdw34BTHCnWWIiNj2tJuQaTuoBTmW
Z2UYVJy18NTXsY2HQjKPRxAChjiDRuxlGqoiSRqN55CVEkW77yUq8tiqvold0Eg8
8dNhxR96bmHDI2tdBvUF27vsffFA8OarCu3dnJYHWvLh2/aY5KoQUpcR60qGM0ts
Y1bgoBrO+/EB3qJBNXnL2sLHQ1Gd7sVDU8HKdOLlu4BGYJ3Cm047BhtDNixQ6md8
Q+YNoo32ZiYUvAdLstIlGIFjsQEq3D9SnghS3pilmjXnkP3S35VwBpH4j871/GbU
f3LmW+Mt3z29wVeLu3Mrgv/aoSb+gYzwNDwtETcnO510WmEJ/Zo4IpDxfa1q7d+J
Wt/QXnNawHs3fQOPrpJOCtANFqRSCU4nc5XtLCENgy430AybmT3ehoa3PRwOxdrN
eJqVX0qsIcyn/gTEO2i45yzKI0nBIg7iiQlK/VXMiaHxUFrtVtcCQgch+GV5Z2Ny
EguGzhCBc00Eyk7kYDXmlpgqfP6IxZM9PddcgXL+VjsYnGBdaczOyu1dsofYuLHe
KhmW2WTTAxqgYaQe2hP+7zqQx8rhq1CMTJ4X8rMW48gH278ci/Cw/HRVeyDKqpxp
vyuaob/f7oJ2FkqrxGe9J6p/I5f0kTrcl6PVt4jCrKGEFMNRKhIpbsA56F6N3NS/
Z4oNi7xPdD6d0FadjG3IG+xGIRYhgskfRNytZdA2AXJzYZLq0eg/eju5gKgNKAb1
lElQ45J4TReSSy+ecgGe29+4hVicuVWnCyarO0qJA1fxfdzcrnlnOdil1fxsFwLE
NUzR4fUEK+lhJo3d12DdEVcw1nXD9vsNHl+AMCb7NpxZclYmbxW2PLtGR/8Uh6n6
pZZtz5a0F34rA9QFRrfez8mj+tsgD+2S1dNXFWcldrLubxsMses7NuaGkVd7du+R
EJNRO8ltzGmwenXifIRJlr3HgHrW9Yvol/T7oxBoC+IlPX0gPiVQMht5rNDP1/Bk
aY8PwsBX9qs60LgcXn12YBYgZxm+kuJYc6SAPZW+FB0xGgTAi5XZKqc6SYKxhSJF
VxH+U5nV4GslcqXxbu2LSgMp/G//xlMb26Z3vngC3TqEdqPqQav9mx2B0kzufOwD
YO9BY/0YJFW2gEluU0YlSm/xJJMn82GRRmB7zJkAP7ssyL1dKx4mNjPjd+3iKvUa
dv3qs6jG6d5hhYaa2/6D9IxpfCXAPebH93VMUhq38chMaU2+CKUQyEU7RAz5EpJH
WNMR7blbvnKSOMGgwXgD38PtBSZmcBe/bJ0VJphLifmGJ5NBCnaB10QpFvSvsGNg
QuUrQptGCrBl6dUyae8s0JR8dEv98BquAVDPsQ1m5CP17o7MlYgndrViPeAhAHh3
1jjZ5w09/muORoMRyUUf7z8BsFgxOZVdvqghwJWTuPD4S9Cq8b1kviinIMLcrCpz
8iXsnMBIQDpkI4qUYO5PK6/vS3hUlXKtJ+Uhvmmc3kBB+jABtwBeOgsQf8F0DGCE
yM0Bk10kA+oWfNEPGu2AfD65yDl7C9ARqYDjVesHzuplAZRKnlIlzbOMIUH2FkdO
m8zTqyToez1Wl7xI470RDkTfsQfbMZGV6GyWEr2Cx3WHcNuouTAp84ZBvzIH93kJ
CBCbqPEh+b1hBS2bJoxxaeFexzbpN6aq93L775ulUNZQOY8SGJu5DpQ2msrxF76A
7luT1hFjGIWNyzjNO8BlWdNw0TIXRnVmr9fUsD1fhazEIu++a2HMv0+cV7XX9qKz
JU84T5etLn1r+POKZlrgLd/niuGAzNb5viLVjNf35qFIa14K5K1j1ePcDbz0AXRX
SXcTCXenbBd3jTqqzPOzXlxg+C6Xj4/VnlsESiK9TAzwQHErNMgUGmTuRCTcWLlz
CCwOjYezKcTNf7b/fjz89GlarsEW0QNFZIxROhtwlEhWq9GPgfmk/YgrAp/jbfte
9XtMZmiaBEwD6cKnPWqNFPD3YfdLe57L9lqQlNaGIMtY96liQPGxFw+cYaFKd+8Z
uKpgUYzp3eyI/BzHdI1UOLStLnLKZ+Nc5AFZrOyg4yOapMDvEMXrRwt/kETyxvi1
F7UVfObKE8cZBkwMSZPVI8ApLjXilLIV1/cTjJVF4us6/k/LrOH9brJorU13kdXr
Bl357qa34i2ieRENZYrRKIOpbsyce1NcPqR9uOtqKttkZ9+w0JHucLC5pYGf/io6
GNwjMQdIjbN053cRouHJ+j9J/cl/GmT0G7noQpWNEuH778b98D7gGayHhSs/k6/3
U2e5yaJHpTTCz2ZDIHn6RrkJzbSUF8FPHJfBJYbCR6Vd4eobxVuA9o2dVstM5BXq
9OtBs5mNXc3T8uGrK6CA3K7KHplxK2tQxhBNILW1Q2VXChOCrsuqW8LKUrh7am2W
81ub7d0mvwY02JkJS2TiSwoYtHSt7a+DR8Es5B3vZ63tOYwfWKuIIe1tpZc3ptOE
1WxomVtwPkvC//HPxT4eD74euvwK+RmgDZYE/83qLPtV+1L0yY7XrNxW3AiP5ITE
0cGiMiVf3mU/c/RiPJFIPOLdjQSdR+YMZ5PLSIRPUmidolMYUKZ3mYDEeaCdJNLx
1eJ0Kjbm3dwLOa+N/F9Lp0fY4epkXcRZrtVDwTg2rEp8GTPORkvy1oK1TmXkT1/U
1MNuIYklKsZ0iWZpQM9FjWhm+dXu65uuWE3LhwIQFn9ne5ZkaJH6UA4ox9L0HgqP
Vpod1dB5i8LdTCDh/gCDmg7QR4O0heOIeocyzAagNGOURNF/xG0Ce0TVPWWzIoOt
VzoIqwiYVY3eUL4Vz1Gc4yLTyAKL+E3o6I7TDWfRsSp2EAx44o2byoBC5vdMdTim
T0RL0QY8mJnZpaK3oEhriQeOr5eNNDAFNAiq5+W4Lsf+V+iYeurutzrNnswN1SDp
xQFIYc2mJ0UzpZd9sXNFdg9HFbgKVfi2pUWeXpMJP0wMlIDYEBJSgRBG1wpufTIp
2HEr75tIV2qnOEGqapyiMmBVpCxORGuvEblxVtQy7MJCQdtCKXyY3Ln2aNYFyVoE
OA/tAezoIDE5EqwOmzU8UeMw0g7HJ0xNLYleR4fuxTsiaLlgsEwxsZfA4rX4ReKq
S78MAqw+yCE/0djlTyMLr91+xfALdVbV4QVtqSgWLdmqm7FWk5Srgxok9bQgfmuH
cnKSqlLkwiyt9sw7zZFYmBdTDadfL+pBfw0nGfZ3Ef3CYHo4KFtBH5MFFzQ7bWUb
+8QcgniY1EaeemmOP9tUh8zs3vmO/Uw3Zb18XP4VF+sN2lCla3L7bIo98X8fDfkd
5UP3wPApffeEgeuRSf9iNHPK0O0YFh+BleOl5C6F6lpQijIuJ+OehAlsBfKqk3DY
H73WBjNziKJ9U4gjpdQUlS8Ny9ZgmRH59j5hRPjq19kwPISwupHbwdpB0QspFqxj
GgkMVXAIoFkjI0Rgvpr9d6DhBdkJjc20cSSlUVmveVUnl7KCtNsQaZBYzIJuHskE
FegbJYyhNAbQhVfQxPzVsoANSEZxyUrsNPaRxuxHTc0dA1ToWXgoH66Ys0Bu2QKj
9r9mkXZPej/czS/wY1s/GrbvI5fpgI0AysPtXPUUbDjReLfNDIK2JKrCzsWb3/ut
qRPZF0+5qWjGiPtrNtZ5ZDX11/U+579KI3UELNS7WZ7eNLSJXe86CpJyTUGL9k9u
`pragma protect end_protected
