// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Ix0tn1qJ+2ZjVuGkH8Uk+QFd3yO11CxvoSqZZWU/mQF19oOwUba4KYJEhBuzvgurS2NNKFsKihUT
ot5/CNeGh9FUvIRkKH3M3twkf/94iVBhJ9KLT7Tn1nLiXm5qa67OKsAxtVIPSQ8pq005gKnHLPEc
mEfRFRcsBuG4+armX50F3aXoWbSR9d6mo29vxAgMnDRL8YdmcE2rz1Q4+Bzb37jcjFQc50xyGo3L
EjPx1Vt1KYd6Cj4VldCi2FsMpEjo0FfVvnVAyMGychUMGSHczIiaiyBocDGJiWlGeQtt2zni6YbG
cuZCxunyG1pWX+KdAJ2AD7MLiFc0tcGjOt9lvw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
MGJdG4BTeXVBc0sEc1gHlS8mHFuhPMcPsvzYFz148FTw3ghOm7zlj9be5poF6LKua5hjqGgnmBrN
GW07w6+xMLwn8Ed0A6otN6p49EKvmcZQxIdpZxTEcZ4JC9bnpWUsxe2DAZIAnQ6G6ibk93zCYJgU
xGVj3RC1WuVjgNSWcHerhtzxy1HSdBNWLBaOhYeg+kYyAaVHp8sdYxWotCLQ+84dn4xvlIlXwfpa
ATLUZq4IRg7Ep6bTgS6xKhlmjuJCfulJd9rdTI9iTT2vbnSvonk9Pm73WvyvME6oQ5I90BJeA6ki
X2J5caZwEEPKomd8GFCTT0l8YH7inuyUueHOsQHHKFfSqF0YiTAF3Jm/pCxiari5IVYQNnuMn9tW
14f7poHagcWsAiZkr0AxA65D1xujlvpvVS7ehkFSrEOLwoV6kjFm0Gf4XbtchAfUMht5R+EQfJek
08Zlp1H+AV9T/8SUgy7GAosRunT4vK4qo+09828jAl0nf1CUOadu5YQtejhlrGqVEz7ZsvXBOTiz
Km+E0svf6a7QdkxMbf6dPGRaT/48++S/S87SRpCqhepXgsuCrI7sBXetW7lRLK9bJsPCYemIyVtv
pTM3bttgs8w9NVdUuuGCZ73mxuG8xvsdoHBjIpTyYhMxqYI34F0YNszB14lYkr2O8Yu61QcARZzz
9HxgQSfRAMGPRyiS1+Hch0f+ISxNkBVevBQnQsN4OFoGfgGL9/fH00zaR+SHG+mcFseUzkMhmTcR
y9I7ig6Sn3tPMNi1U7LgMvdJHf1qdRmu/GtskQ4iTODkUGBCbSOHY4hxbZV2RdOBHShymV3+f+jE
W9q0b1ibdwBMBdVnsMtHmhn7Tng4+WwDgifJTfdoQ2X8RgZW2Cd4VCn3Bu1bmC/PPK+j0PmbO2Uo
PFpkAPOKxnxuZAYvSqdc/NJN9540nYDQtU01qtbhGbflhhFmBQPXr8eG4f9yquLFGEvIev0oFAAh
kPMVOnxItkDptgVf57O/2IJ4nnOYsaAxiaCc8rvqbsNtkWw3/IHrBEfzodpG9XjonH8YS/vYyXum
K2s5nm51O1QZOEj9wgm927BM/qcBivZR5nnKwGFmyoTCyyDvXM59Q4VIN6JL+2/8/TfIZqDHMNLV
ieFt5CBfmj1T7i+L/TOjb8rjX0AHhY9x2QCVcYbRPn4LVJah5spyuGlpCU/HwR4EY7lngFlUIxsk
XiGQ6ej2UurO7cILPz8rltUq+9NLgAcMNkicaXgXk42GyfS0FEOetdu/QOEO6Ut5dVRAsGjiWiMH
Dcmw5Qmc/1dIpZM87/zMbZ8ZfpNicNtSIfBy+dYCBad8uOapB80WOxv1brSII6OMvKN5EaHw0Opz
OSP5V7slBwzzAYSOMHKORiIokZp7dMcEr/uX8QBMYdodHKTYUBH5bzHnIoGFq3uWm3jkcOCQ+2P5
t5L1dHITbg+o40N4vzvXhAE8lAqnsNCaN/EHsZ2nD8Yy4VIIW+iGWf02PtBsETycEUc5G95mzvFb
mE88dpWjcZlAHKsqI0G8zT9kNhKH+j+1diQfETBErEpn4qaGMUk3cVeWxgyDITAiYLIr4fgfRVGk
OaifLQZoWUCVovym0dH5awMbeuS2U7M30/gQggJX8L+e6DqCDjPronoi9XqSYU+9c/QOuhouMVsr
EvGYz4+ivW7O4QY0mJUeSHQTyvH8VPH1qjWZp+HxrkqIwx20SJTGHKVlGyQRx10oKKV/LCul4rsZ
9bfNlzwkG0rVhjRnY2yJf8sypAVUVvd5kC4LDz7xiqL4bgShdn+1oyMXPDvKMss8vNpan95v43FN
yQSWiRK0le6OKxVKz84l2C7etrInhFDfkKd8314gWxYRseOjtsQRmSxKff8nye4JKbjzflL7nYOT
T3k35fAebJoP1zHcJxzpvS65rjbunD961i/pAedzHdJTlf7rYYTsHorPOgp9QQ0TcHiRJCZDF+l/
UuyG449viHUmESzfHVbffBNpqpOJS+3QQj4zWDRuH9cizIjhIXpn3ydz247SIYNBCSCnIHcXIPJX
3uxsBCBhW2Q6D/vV5DovT1tSHxXt4FKK4xCl2s/voXRRdxSrlHKmwWP4SDEjjA+DCkluqkYWykpZ
/OX6RuLsHloZpCe0jWS6XXzsMdG1GZAQ3+4MKb6iLvgSeYEE9tlYte9X9HtI32ZomdRdW51ocBTT
BExRmpax/x85bu9n4n+vmQMVWxvtnDVbsLEZdjrRqiWW6Dqr4NbZsK7Ad/Hu5zZNn0koDNP/OE6h
t7pD+gLyOyxuHl9lg0ECcKBbARRxzkgBo3ELOMohDd3kpNYABi23UVWZWFibtmqBcYwiZ0kS9hH/
NU+NkCAIfl9UA63R05VpfFdb1JAcvyWpIp06PmeUTj6gNRWmffwfBsyVGXfMW/IYXC0wN0dwHcP6
WgKZtD66l+Rzx0uoHAm0ToBIjhYJoLpYc7+O8w9wLpPpLgf25Z74ajK3ezpGinIG34LYFB6V0LMa
uUPxhCW2YZBitoB/BMzCBG2v3l9wLbhRxqSlQ6DxOpG41M697WwnQwA0LE60zpkTIGwbJeZq11Fm
WtvBvlg0aSKr4ZmlHcE7aLutXg6m9vZ4pzpIUtVzRw+Peg/Uk6CtXQXH4pzCdX6XMnE8DqEiZX94
Hgor2iQkIYmXQ6DdcrlpC9wjkQlsqVznISRK3u+7sDDLt00FGP3NX8geDlKXoBOo9p6yFHLKeHIv
C20k4xIjKnvI9IHLIPv9KbJ1M+9DCFSeGx7rAwGIitc4wiy5ndqvU2YwalWP5LIQQtCx/nHPIXrE
7AZsJ25WzMZpAjTrICDcIuVRFHVFrZ0j9QtPhJSkKnMTFBblSmf4/M3e1fMOIgbEQBnbtP5Y5d86
lcAIrt/Od9VJwiaI3q6/sypf+2dQv+CZN4Oll4ZTagjDLIl5qHT1r97oZmbZ+6XB5ooe2wU6M9VW
WcTN4Z34UW06Yk2D2W+CW88QtwfnuHua96ZqM6CdqqO2wtWAaj/kAmkY+q9aOnoKEoMOs/A59JTZ
cD+NHLS6eptRHwc3pCf6q9z3a6DUnna+DWIUzaAlkpgq/WNL9QiMuyUSYFI6IxEokxu0wFEzfKL9
+6BqAYWnk0breXvTHDzTktZZSCoyfIKoezU70XGS/adMjSPhefpVZQL81n0/npufEu5fJhDgchS+
0Ion0ZJ+yW19ySRsJ2Bl85END5V72JT4Yp7isGOwOjR6M6svFuZovf/nxr4udqitHo7emMeX706B
uvmTEF12UEZ2HbzHxdYJ8mlRhPrSzXVBnGkIOiM9jdUuvWqFBt8MUP835tNdPXr+mtMfIOPR0UPi
or9p+1I8ZEOj6S6oXDEUtHiBBmzJ2czTO+9jd2HNngSDxn3wUXuPhbQ/BnTQ79MletEs7L+gCfn5
AUODnfrvrtje6pDDA70Vv1Aysq6dIRYcYuInjTsHHA9N4P/8cLx8HlJsRYaHdtkZLWyiutMCIr/O
prazrvRMPtUKc0bn+WMY4dqBpRGQ/5mUn3NqPZshYFuHpTFtB16PFmkY/GqbywN7UXBfg1CcjwPV
6AdtexL0+7vwwEuzOVkHF/S2usYlpdAeE90Dk3/7NhZ1hBGcZHM4MNvrFRlSsUVBfYiZs0fhjkHZ
qLtgri0DJsKfsG2NaMnogn/hWjNKrNHKB5xXEXQXwtRZTrw3ke5TA0FUMt7x9OfWV0fFkXVoGOcm
rWK0gODG8OeO7dHPyghsxwwY6r5eXE4zjpT6yH6hKaKn7fglk4zKjJ6i0JavicmDG/UHJ8QgVuTG
ZKC5eBRHjRAXAQQwqnN1/SvcZLvZn65SwgAbXSzJbD6UrBHkh63/M2MXCEMSfOCrM42djnIsKtFa
twkImyz2NuEBbpAoI/B5JVelb6t8u+Ea4zrIvG6s6njkGhnRZRa09VHwXQGdlwU3v21/cFv8YsWC
9fNMnMW8em8RxOBQKBET/jqunS/udDEpU3zAKJoOoxOi1DfgDCr+7ycg1//CqwNYvUuwkzJdc6NL
dfenLLSMpBtIAS9CFqooOyObGpDaeRK+IfwJN8YJHnaP2ahqGQSOTNYTMfg8zSloFNpkYcEpRhph
myBm9VLVoGMkF+WpiPU9NNx2WoHJrJAnk7u3kOi6EAQtdCY3KJ+aKx/7/SM5ikYbOqbneXmsjjz3
M+RomBauc800s0FI7KqsRfUDv0sGI7Js1DVP02I3E7uZX096aCJUWoVCcuVNL7m7h0Xn0ouzBW+7
rbJa+TtiATw4rJPe05pTV8NQIAaZ5C5oXwT/LBI2a2+GScAt45/hAHKuygf/NPapZK9vMpaoAJk4
M9NlYW8sbJkpAve/FneTTswo69v38R68QOaRBzRjPjWwQ180JhKAcV5zbLkpvCNwQy0C15wUwQS+
t3kDuxQMPkV3FxIS1vlrBtfXPlLscJ15CTHa4e83O0eM+lOEniTPg+H2l9WggXA08AsgtBK1cn41
ZiAs95Ptp8bIF/qlkLRKEnu6zXIanMCGCJOyhXajFXQs/QSIBCR6JruxJrglVw2S6P3jHAo7Bust
2/iPwNw4em4p3a3a06u+i8dNnxvEzMHFFKJk9goGCqaXrWFaTxFwF2rPFZ6TsJF7iwfTKc+GG/Ho
zeBLUkX9YvTvBrxjE+f6pGmJliDj0TdndTa3zFPpYIlzi1Upqys1Fy4k6digUfXe/DVZwn1fcB/f
FOLFXNznxv2mUCeqgrtc4AhBRaRrpipKwJKY2HbSrIWdVXSU7Q5iatsH6OXqQ1xpvR5VhINMIeYr
rduISvUzD2F8slWLCN1bIw2xDgI0DXGqa1clkByLP/OW08LR9uEVIm6T/Y80U3ihIIbxXEgZpHGQ
Uzio76ELzwUiHBKxg81ZF2vFqLSEwxkonK3tFt5GrpJv1mfyzvcEbNEIJizQMiA/9UwK0EU5X09w
KBWYGlDIQ8wU8C/4i2MmYgvP86NI0F7V4yuBQBLlGIfC5dSouSfPOceltQdt7d39ZV7xbTQ6bdB6
7TxaJKckAlJ8LQYKFCHmReOK3FmfAFYSRW6sUZFmUevXe57V6ZMCwemb7XqQEB+1x7DrGmWxQuoO
4zqTLkUHgoGIIW3EjbUSSThzaRGr1oWDacB7IKfIRig5q9Y7cBITcVjohhFDWM2/X9MK8reKRIqC
y4RKvp9/pPBEHAWONGu85vxsT0b4S3sBostMK9n3qZ4+YM/n0uWAnQezyADgFS2ccMrwsiu1Jvcw
QqZW0VJJkoozdZvndn+u4zkyyK+SnXTddDWkTne6POpM3Mp/3Ehqa0t5BnH6Luytxl5gAvq2nU2C
EdiBtHkqKQpGsGnlLZs0QLnyTJg64piht0cgBx6ssHpvWfy4shz67LYatdHfYJOvwBrAoUe2v96y
zPgnLyZYNiFBwKxoEmjWKXih3lAo07YxRnUsyG/Lp+u8mADp+IFa3m6QmrZ0rmXULPPWlGWESogH
IXnR/r8yL+X15KusX4kiGZOfgX9Hd5BQz9HWyFKz2OErYfyJhh5bpH4TToZtYS4/R9CSMGXjPDSw
G3q/gInxXPISfw63YqtWwy0ajRMTfQFr0q76h6APKVABgfSTNPOsYhpZe1RCZLtXcubYIYdiGRlx
5iTZNBxQ7T0vSTL+PnoYlTF1J0YHLbEWI2wX5F81il04OG8Ujec9hvMpU+WAGg5U0l8C2nyU0ccf
Zzj3Myp0fpjVqqk0YmfCM97ay6QTuJXgJXa+xW/lPvIT4nWQWJO2hzrFNpYRBOYMO2UuFqfJ0RCX
I9ftiJ1u03xuNVOqt7aeACYM7KrXVqQPbJW6iozmjgOjUVnGSsTtoQ661tRQ0hmWadAiYYnCkAV7
YVS3VlGOgO7I/4V/YRewK5WlV2dI5KHp95U3eZAYzxYNi7NuKGcq0Js2Ey/W6be8bmZtUfO0jY7X
dQdQ2N4uT0x35N0SzUnA7BBYZGOG5CaGwjjCNMDcFI2YYUVjAJoDjR+n7uMwu0T3EmEYv8UkdosW
A8NH6zScP7n3OB6JP9qQKS7cl4wNEGxLRzggxIASsJO0UbC3I4alh+BZhwSNxRY454mZb4plF5mD
qwMFlRPyibjdufXMGvkRD2xnE14dgDikSadWd6DwGuC+1Asq/SKftxnfBbdwCS2cY+Uej2I5jqWx
hk/Oq1nK/0PtBdMbwAVLOQIPhHl2JQYAuTKm+BgygOZ2gY+azGaUXuIwzurCdNbaHaDR7c42zRO+
ze6nzquJI7+L+7CR+7T8VZG83JH5FU341gllOQIeYFl5MtFxbGIHLDS0zVhK5ORHQAtIAU0t60se
NE+N9NRg/FNpTe8cksEhVWZFtsE71C8zLOt+RTWqPbqsKZI5wm9sdGxqDgRCKI5tXF+GnVlOznjq
I8bMVX7nzwFdxGPD57W5DeQU9KgmJ5zWPo0yOGMv4VILu4ggFCVUtyoUr8Ji0cSLzJlAeSeJqg9g
37RSTxGBQUdWX1a/J5c0HPA7Amuk0QTiDvGnAtL53YErQfwcxlcELkhEPYWJnbu7nu55+AMqDPVr
yWVHGjrvFpcVyvHctgHTgF+b3U+lp2YnVP8VqS8EoAXZYvg9Gt2xDugM4DQCT5mdUzfjbrPoF8Tn
NuM99tU6BypFo1onYANR6dCUjAR7JCiBS5OYaltdUMNhakU+ZlG+9tNsPEYWGNL+k33Kq/YMiP5e
80SsJUgpIV+/eTJO/grLxc+E59Py4tY5MSWJijPF4rS8VyZ+8EdXDIM5TKSZCN73TAPjMxYNzVlR
qBy+Oe3sbdqiZJghbYFwk5RnlG4CNpiHQKI5pZbFns0BQWppoAai60J+b2/OD4qpAhramiSrAoiu
SlbrRsyshdwShDsZ/H1VLnkCg7hc9R6kghYyCAF93PFBuixL026cFwV3rSVPs5yfBHnHlO1oy2LX
kDyk/V6wZAonfFgJNL1oaLfFVGddpmbg85VHVgl2qVpfMVF0iQJ4tekkHv/yCeutZ1PLYIGLAgoc
s25/psrGEDYr7+OIHLHVjdfFRFPQxqkE4IFMlLSvCVOoSoQA5Mnr8Eui1aFGTXzyRFb1bb/3v18A
FPyuqWEnI/FrAdiW/b2HsK1vkbD43PsKE8iCVgHG2A4XqnI+IG5gjX8fzv1KPjumrZ2hfZMLSEo5
eiWk0M+g8ZjyJP9WHfkPA1LlNeD1CDREdROYENV0vg15ws7f8RDrwFSNbZkMsVH+hRDSRW+SgCb8
sGEaAZsg0YkjRGO9vrCRn5e9cURz0KSTt9JaDELtGkeH4JAHA84aPBm147ROKXXy0J6K4zfh/1Mx
UJyNUMPBYPZ2APtwNmFyuRxPXWKoNOi11ny6Yg0WpKMcc4cREbEmVTzaciLjvnbw3CU5E1XDuptC
oBLlWPbOHJFVoCPQxEZLBQHrlvuZWb5o/blOBpM51hKIFQvQOI705Ba117B/AxjdmBfq45pWT9NO
wxGzeTnUSqN1Vh5clG5iAys2p6pqr0ZswkGAz029beuH0yWJF+L0lLUsaRLG87sKFbMFVx72UwB+
sIF9TkDNtO1f95qGQMoqZ0gPKcQy2XNHLoYcZJugqUbJqAbnRxVIF7cXFIp1JcKfLTxeuQLV3G7d
fjLLcCuZFEDhaQyNQ42BtDSLmFupW82CM4W+tHHpf6C0ajXqY0QHgO2qiXx1fN9wtr+y1i33cLXP
BEb84lyYUyO5LB12ohyTY63Q7E4FsjnzBWfDefyo8+TVrUXqVnBNXcw6sufb8IJCHguIQkgaYPUq
X/rEDBizJPWM0cvk99r5bbfOcVsWwpDrYQbOt4q1rIyj9rysm3GfzhL13iNMa+ypaxqI/VibsGZM
bsMZPKRKJUl41zILf3xUj69Ael/dc6ZTch6aHUy2hJOv7jZTC9UnTbaZCvdGUjYE8Gjjr1UvrIJR
JsKu29CHTg1A3FEfij0buCONf21ZZqVam5vAbHXCK2kAYeVt87u0p/IGZxefBk+I4NGxcOLtLd8F
x2X+vpiTv6ViBRE8Pm62g6Ch+YRRts1ffyO4eHatPwkgpE11pQJQ8X5SN+l8ypzUwkolvUzBbQfU
vup6/1XJijQheWTJtoZaRNa9+WMk5pn/KW1a+b238YP3zeNOnuyoWLqgqvGsZulg/O5/UHTQDlaX
fx5sBKo+7HJYaBoO0+qUrudFuhR9inrvSV58IfKks54XRtq/eBVz+J7WAz7Zo0EGaO3v0PfDqTNq
jT106XFJ4SS1etfPx0WfTpYxgLMAi8UkuhTeI9rNyMvmVv4ZeQf3tvltCNsh3A1PVIKcDoSRmJfu
4qNT4wIN0uwGk9jVhS/hRZNI1OZlBS5xwfIkWeQTMJdgFe5NSOd+KygJSdSs3JxvAKDOdCMGVzkd
qtwt0RoMl0b7R9pgOX+2qyb3B9etPFGQqfQLOKCYmb1WU6FTNKAMxhZ4zQ9Ar34fAEFSMK9j77QE
2Y+nqU8z9z+UD/IsJu/Y82vf+m3SSzpZxMxJDfYT4Z1NV22txN/ik02NJhOVh9S6wK0zy9ptYtfH
sClnRlCumIRjCQw6VDzPiqUybaFbRaxV6mRxjliKwa93ZYr5zJkuk/g7rS9AZH2AgjOWberh8ouu
V90f5hf8OiFkMJqF0BAcybCK5xfZSds7iFlVQNlGnLn9NEV00E/BULuEDmUf6nPKwVfpOyO89l1o
rmHF1SgN1ayO6ES815S54yN5bfqs0TQd2pBAmbj3w9FCTf5KlmPyWfFcNC2NDHAc7fa6oX2dD2Ga
9vupAFdGJbb3nemW8Lma1V8o2CwArcxAhYnlM++9P1IrwbY9VZi+bkq00sfYqHiawiMlZgj7PYw8
xugSikHF0gMISe/eTxLXUGgS/swWdqprwNBgnTx/jGMxhTzdc+NovkaLI0lGxpVqj4iTrbnmsQ8E
OjUNo0sJNazfFEVDZArEN5wPIcykUDOJhVSQJn72f7M6/+xeLu495nXmVoUs7cTaihJQ8J6EHI1b
+Ne1xZJfl6oGzuEMwuO7zwPYef7rMRwIbwyhpD4BGyPO/oYfCKVZE/CbdDAcWjj1qLHkndwWYzce
b1J19apIegP/LwDePpDuvWoE2p3Rz+jyBBgUt2bNaitAAnyBV7SuTNRYJVwIFZyaN+qmpeGUPJKB
unuVWNahgYPxb1Bo7atGpeTUzQwPwNL6IoiAhbnSnO/uO5MWmoY5rylgDNkrxU4QApFdgwqnyZhY
9aXrKhEoNaKAjHbx453gAIpqViSEUzyjboQ6/GN6xCjaW4d+Mc2C4ZYSUlEaEBgnEfULY2yIuZ1m
Q21mrAU8UuhskvpS9Wp5Vek4/bvPjhXSCwNy3UTgolHMkjU+if5Nb2/mfQjKaSMX+a/ppHG8/s3a
E8iKNQDEVrNSfbt/I8GThm95FrYacQXw06E5dougvNDzRORNbOblBRbUZUfJSyzkFvfdZo3/DGms
OAfaddu5O+IZQ0/DGMFu5sxnZPyuGJoQbAaeG0iPt77i2//ZVyehcFZ5ydqi1Vf2kT5SsoC5fyui
rDgavssBh0ZLkmst9ni79PDxq6lRef9z2UK08urvIT1Xzv5B1LxLUEPFpQzIyeXt6tdJtOEo2wdJ
LQb0eun0OKuvC85WD7psgVcYdvmYFccNomy4HXWm62mHlaszXb442seI37xwpWBT0ww2UDWfDvtS
amI8aedKSwyyzNSFkeTslzS2JwlL1IYaDzfI0SqvnjhxIMx48czDf1KbyUK9HmPfuQytQpEKmAus
IWBO2A62AbNxt3iONuI70e1kJMM7EnLu4brrNKx99C87qncboAUIeY/9Pm1APvlsh5ByTv2axv0i
sy0N7fpF+4lFSqcWaLJxFruSCq65+XTzzbENGLc7eDXMwQ9ugGcWPJ37cbiRXrQ6cmzxCnwQ2BVP
fvB/MCB1auqCj/sGOxPerx+58MBCTu5RZDd8qbsVBqhMpZcZrbZf6H37+b5tc4Dgz8ECnpnYzn+2
MwDiHApzGotgIZqwuPMDgzUSYOai6HArClFmpFwnIXgrydaC0agIAZ2VENkE0vK+zbAWAtWxQRYc
7HGQl4bpE0bhfw7cSyAWVVy3tAM7hpmwNr8PuZ6WHmI1hIDKCtEkIom9QqGflix2jLQC7W7AbbC+
bfOdvZCsY7Yee2VzizgFUK8eZ2KHph4I2foG1UjNj9YA91YY6Z754oQnmGU4HZyrMcFXkpCHPIkm
Uzds+SsN/6j3HSeL5Ajf9Mbnq4K4GQMqRJwPLS4AQFg523dv/utbBxIwvjzrX8Ltz+50SWFqkuet
XUuHhjKSt90gzRcgzewXFYh5dY92o0ueE7oVXv/KwrKG0pqo56HKUxRZQdJAvAVEZVPD677Vx9jB
hjaXwSrAAg68ugfbwOEp+kO6HtoI/nhN5YW6VE4x286Mpik56xFRJN2yPs5r2k/jz7oDoU0G7OUz
7hWgjuPOZ7ufK9eHCskrjJdHLQSkk4oE8WtRPfLfUMyt29p1WaxwgymhdQHbTektbvHxcOvJ08wL
yh5WqeD+9MB5W3XfrerEoediCpaQ3piv6NLDi7j48l987BINPCcPCQR5TCcV3wqfLw89c1ZaSmjU
S6HTdI67qj+YGzRgGEICGqJk8DmPOYeaTF80nzsrXAEOTuliQiGIOD3GU6qdJUuFwSYmLcbdrq8g
rjBXt8bB1Y23L6QWsAHdljf2EsTxkAC1/K3P5KUbwHm1xt3xPH0xaEfqhH/eUczJTJjagDWynwdv
IK2o7UPKQKLGHsI2udk4qCnqxAJAF+znTT1GY3qynbvs5v9TJC80kg59aEcLnWzXe6FfAUyHIA/o
RDAqNgq72Gi8ZNK2TlEGV8gtt68c1p0+mXMrtHeKqz1MdBCCftk+q47WDF0kSLgzLrUxgTML1GPt
7+EcvGD0BSKSuK/ITH6TBxh4sCGKVGf8aUYADL/XbmlpwJoO9jZkdIoXLlv6u0cwgvbZvOyPF0Ko
CGzq5kCK5j+CHV4s+7Q6YfWXr0hNMaU8gV2ew/Fs/KabuEdZsUZS7xDGGqpwT3Z3DKrpeJVOBjFi
C/zC0s1CsfSZnH4JTxxZqPNUHb21DSVMKhpl26HGRbJKFS0UeLxb/+yRVPgIfnCe9uGnZ/OZHW7S
IsWwmx/18n6N3Vun3P1n8LX2Y8Ao6nZ7BYgOw9CVpWNoUDlkZ+5G/zV4YsLOs0tGEnWYO+q37FVe
2rIf0bIbRZUVmL4Cuj5UuupMboix6l1vKS4OGsooiIyl9zLCBY94k54uK8mG5VQC7xXIW/aMxlJN
1p31QuorIWKPbM0H90JKf77B6WtbLjMAx8217eNhKqHKRcsvNrWQDRmZN9EsOF/DR0eHOuvcu1Hm
CdCsyKajSs7CgiZ65I/507V9xoQgPESV+zRMyMRS/3KptcLqj3OuMPOgpAbrPGpQQDYC1LLi9H9l
wpemxs8RTZ7Qyyic3PRHjTHKejITi/7gOvRkFOLTimA/JpIn9tx9x3kIg73IMzr9yNO1LHaIEvAh
G++2u4vcRAwIKIqMyvtpw4K4QPXI6ZEOy2q63Qpctzh3FjzjueN+S1Vtr4s1iIhH3pXD75VhFnEH
HlDFfr9FO/8TUW2DmWOvl/ZFbSXfDHy3raCcKgjlBCcc0a/6do4V12WO8WrcjmIGBoOHSREOM2CH
/3v/+hCqtT3qEkIq2IitOWmZsAJthdAyC9l8jSp4Zlz929hUbPsVy27brzCAmmp3dtJCp45ENFTi
YeplTD8hiay9YHECQZtXwjaJqxcAOeKjWu27/ZRc4GJS3SBTgtL0N1RahGpynIXOP/bckBwcW+0E
b/Fxrm5Sdxm+4Dcof9rkTbF7zG2N9s2h5Gs+WsCbctgga9eYOHqKC4W0DKyDbnnY9L/dAdmwEFQu
mdk535dITqcJtr4Ck+oJqEIbqE8euMZ09e3bWMuDMB8LuPXQQS4zvwZcsAz9svXqduZL9H8u6Kww
ggUKDvY7dcxeJauNPg9kGMv065MHofqf4aLyN32SZAoDIpmlf1vJRQwaEXmY7oaGAOtFd42LRw94
92irKkBOYhwuU0gNpMuB1One+uffUcpr8Enrxp2c43hy+a4CFkoZpZTr9XkiJRQEPsRYeMkSbxyo
sqBZEZrJ8zNHCZFPxLy4YETn3+fgPAg49irs2OJrmHIRoyIJLykYj48du4GvqdUWGXcck8TX2LwH
EWCnUXTRIauS75p7qlnRNgfE1bR4GBLTkEUvBsrwp29WJ6PMVe1zx2z2uTMJTsNoaE8021wBUUBA
Upbni+yPi5du+BOkBO68a9cRX18mxN29OC0K87D5eeD5XZ9qnExcEv5cgB7w2UtgnqdnWqQRHKQM
YBgEwkCasBa11ZrGoeihvHZQJGfpO2tGfdakoLw73FpX12NOOkBKQqHrNcUJr2w4pkIRenJHkH2j
66h5EVXE43FdD8KPiOyC8gz383EivA53iEKc6ShSYBIM5nqTTltDaShtHiOqwcsGWNzPsEs02mVl
gunH84IMdOF2SUuupL7U/OTt6uR3jpvwCYu5E5JtF+a1iHhIEGUWc8I/TrZhQDCMWXg9cnZ8NtkN
X0bRolZMZme8UQMBac9ZHgU1BstDMvbpn6awZZhRfAQqKjpdXolaB6GZCsJPXSxkmSll9CrRrt7F
UDK41p0j9EhgJ0dLFbO+EZMiLLr2EimtaF87CofSsMbVMzDVdHNWUmWZ09iYE1I3Of8Pkm56bH8P
sSAlgvA+//rz/f9YRSLQ2iOaFqQLUDgTMXMB3C7vNofG6dniW58z6g/hKcv39W5tkhla5kOsd3Ol
j608YjpIQe108UVF8FNcZyB6r0bVf9H05Ts1NrYVXrk2CoFXWh+0Obuzbeor9R6qy4fBohzSdzld
azimJcDO94BMtauL2gKGYu2HlG3KXLIEjYo1LzHnShiAjXiqysJ5GWd77OP9dzk4fYX36dOVrOHY
d36JRpm+Du4uT9z+qG5Dy+V++3tjrNLDpJ++zdkOHyLBZGAKybGvGDq9tZlzbdaSjRGo2uLBztek
mHK+J1aftKgInk0nIIHYijyuDlZdeqRtepeenUbxtWEnq78AP0db9e8+et2yyD6oJ8FYcOwQPoRp
FNqaj8SMeiG/AnjTjxB6wT8x6mG933fQF1w7QPO4Eg7p7ndh6rxvZVeASFZq0BbDS/P5I8oPdhQ6
UTjlE2T41ZOSGTX0eZtgQQsd/bHD2R7nYKfO/Srr5bGz4TZjTgHqxdgHvkuyJ53Hw9i66+X02aLE
6NP6sq5MTgPCPb97WwduvOguHS/9iI4o09wA8H8Rkd+c6LFiWQu3Ekp5e7Wd8XL8/Hot/kba4yA3
xueVFWEQaevasNctfz+vlP/7Favb5gUg02whrMe0tUN9OYcPPWl5X+m681YL+umAJmPo0UbhWwA6
SF21VhE8ODmrPN6zSz6kzfox+egJo4L/GX+aZsz+30a158tFYs0UkBWzcIHbHy+6OWc9GloFsmb2
C/DA0YiURYwkg14RigoLdNN97Py307YDm421IQKfPUntzbwWfQ/oPydTbeMe2WySr2BOJPsepkO8
lv1nGWUVsyeOWnqkHgai9cj2xw6FUpBmdYyWK85Jy1bUjK3QBzoIk5il4qlhu0JglIy7NeMN+n/P
/imcJNs6onAeC+pvmKh41CuVDckzPoA0HLyH/bpqqnI8hLXK+LP8EtW+RMhqZxdRsKrFW1Twfe2Z
B2uzeVkDBLQVSZeqyVrUUjUGRJn1VkkQWDoWHK0HCSxkJ1VihSXsfBvZe6g5UkcVZkVa1kXLTUjS
PT2XURzakR8tswVtLXC50PdjTCn3ltsJ/F31rtN42Yd4150vkZIrftxUneRRQPjwhp7nCApjb2vH
WhXKdZMfONtRi0D4qoBm2eAIfkHuHkYCbo6ZMxgAUP9ftbdFQk7R1WO977mbhJ9OyJLzAEIIOcro
XgNEaXFuEwC/wx0/uR+kAOWF63OFHVEmyGSab0XtS9ET/56QnSGOYlvKW4dkJlNwG/sX7WkqeMLn
14zLbQP4qJ0lnFtMWw7sO74APbiWs81vKSD1Xvtk+Uyjg0wVfA5DSxjjHYIJpvmh0v/jqVEsZsQY
ydw9isgkX+VxjSQxf44475RSB2u3FxLn2/Hs/8wYLiwO5Vwvx1hWPOiFwK7ts4IRU+Qb38vVCpPd
nbTwU2NqOWFqtbJ/UdekPLpcRLL9mKbFQCyTR0nfeYiGkYku5RDWB9cQNo49uun3JdMdhP0bGigw
kZtLMzFGV3VDtPbOgdehaerYap4jDK0w9kVxIbOfLegfIt71FAuHH6Wo9jMQ/gzdnl4TSkBq4iPk
cTsgIpIDx8f7Kf9oIEMcJV+GCZjuJmxydncfgFarsmzug+3vAuqQGDtRLbKhlVH0kmDaFHdNtxNg
P4Fn7sU/mB4PSYy2nSg33QGgH6OeX87jc1Ier1XboG9vZicBzBjAAmkV4s2l0V6aGwDiTPuC95MZ
SdCWYzcbiHMFszjFvS0cb61F1izWOCvCgUnGaHHtkhHnMfkZ8MgnbbIdgpguwOZcq0T9gqL+aLGL
J/KH+g97DV+spMU67Jc8OYKmxwYlNn8Na4Te1dgEkrfoHIMoDFUtqOZ1TArL7XmF1t/Nz2MLTQe2
B4Uzutd145OmGZXlG6N+Ux5iBqGortGQwEPU6p5tL1ljrQgDE8UQfFP1vR5WiDU1PZJXcyC/ReSl
P039v/tgTH752oNrWIceJqf1KX9lJX2Z5QIansmIbq2B9Wbh2DM3VBEdIZya0ictUSFlB+DZYe6W
UAO3iwbO4QZIkx2C+ug1CSS9fCXLExQTmGePaVcbgaceNm5b9DoXf1WTIrvPp4dtAD7PBWFw2TnX
v1JAP6eh/gcpG3eQdgdBAjLJfLNGHgHf1XsMZVdGCKRaq3KI3JA6usN4ldO/9j7mBxSnzE3hsBmh
igm0p/x7ijWJhGKM273px0kyavOzBEcJm/EYcMuzV5tCY2FGXHa8USbnqM9T6NPVDqClLjNJZPUr
n3P145KWBiUd3yjUcpRart4L+YeImr/7Gex4IkQzWfLEJbtwPJumIp0Vi4CRW2inHlKjXMrX/hZ/
wY/KQQZMoq38clgxdOGP98Bqd9F24ZlMS8bf7aoN18p13jwIQ2zftgn7KuJ2/3dsOqglm/OFtDLy
8XLTwslHunc691pGpt91Wnrajpp8igW0unkUQ2CGZz/LDWay9MJ892yIx3a5SwgykOP8RHuCJSkt
FJqyR+q9/Z4gTgTXHNBmTskv+Rh1Jrtc/FgYVTwIA/s4PDoIZey7iXA1uaQR5hnw2S2YSQ6/WzNX
ur1mPcUY4WvvGP48Yq9pykmGWmf1mTQnKjLx6v5cDWc6guwXdl0jm0w3IBUlvXp0M/lW+DrvYdVO
+FUXrn0dKoVcjqWiMnpacuxwiqdTKHrjQ0HBdiYoeEU7/2zBPcca0W4kHIKTjNszFl6c2Rnk3pB4
p7P5JPjOFj86TbYUhiOsQnKTQ2td4jwAoKp/RKYqarI+jXIr30g5ZBHZn4Zh+YoXFVTW+VLdU6C6
rHap1JdQr7ckUMma5Kha2UxSQW3/Vaobuqbor2QGVZOfK/VZ1hIm5SIAmfbxb2PPTfrW57zlA9nC
WuslCvLxc0zOzwQxEz4KPRrB1QupNFfsHZAQKAUKDuH0YdUC1rGZB4T8kyOOctz8OtO8wgNkENWj
vctrs3Vu9nahazVbPhy6Ur+uRbOyx7a259CJl46ipSbZuSUrDF1LhLl7vx/OAYkBx5jqv00uP2xe
omQonzFoUDVg7o4ZMurK+YTmJCUigELWkYUoYkulrmSFnm0zMtm6M+rDRLKHt/cyXljb/nKIffp7
mRzScsuaZ0Yjhv98rvZcJrQ+QZIS33nE5+wSSAUGmY21QPcbn0nMpnGwQgEJ5Et+DGb0TN77sJRD
AG1Rj5kpR4zFKosbB+c2dBoj6vtk8C31omlpZ6grDUxZlSPhbofhpf49PhbGCVcWdaGf+aeC7AJx
WTzUcZHFshJV4sWuK/ZdoiIauU8wMqMMeV6JomqmRDCQfIckHzDcZrJgPT6zyPlLUs94wkGJKrJo
odYFjVuNLUGdlt9a2GZCGnLJTK7iE8Qtz050t5tsBn/S/KCxnDi70nAmgEsHdRxpmrEiE3+hUXq3
OpSFel40IfH9OMm4nVOo4dKUZL3gzPrihJBgeB3GY1e1EeItufGyw4kjZ79h8tjVES36brzQktDQ
CiNwpHC2VJbrn4zC9AggG96aeg==
`pragma protect end_protected
