// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qGnivov+In/wwglU2c6WMaDANex3hqn6hNj6eZRYVCEvOtJW6ihzSciYgHdK6iRvJ+Xu9mRiQa9k
+EEHfO0/pFz4KmcLmycAwDVSZzgWehFvynI3vDW0Bm/nv1OzQVNzF0k+yjWkjaAs80i7pyGg7gXp
47S5heagVgRffLimDYUT9PjPx+NRSiaiMaUljs3AzbuwkzJXKzuYUcUmel9nGjz8dF6jTQ7rgOjm
ubhfwuVhmcdKbXorJhvV56Hchj5SGT7L5Sq9KZoHIfC56wgATFkSsfGtMNODjztSTAkMkuzUV8bR
MMfMqeTk5NZgWBZvFQjM9NRUkwHoST1MS6jAbg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
wULvKkMCwkc9YMf7ThuRv+qdkNsUCZB3DO/TGTQrGcaEgM0edq/AY5Pfg5Yl/S5hwNxHv6ViU33Y
vE5VE1S5eR2Jz4qujgCi9AEAklmNu4sG1J91ndsCTTqGjBXp6qThWf12xOiOZW7vG7cUeWqsKGEE
+MYGoVkUPi7tOf1KraCYJXjmu6zHq6DDU3YXvKNCVvEwbzeEPEpphVGsgyY/O93dT8GMvS+oxhi1
OiB2xMco6szph20qOkgPlH3In1B9W2iwPE9W5N1fiXsiMeuC9DunSKVDg2C9rhLzFQvt9BiwA038
63q0cJw48Z4Uy9A6FYeCMaEGJSSGAP1QRnPs93Eqf52Kv/1UvZ5UY6SIiZgjC9iQ2JR9IdxqHl4s
ix06fKhLWhfztU+Mq7rHug6y6aMppUu7KwdWa2YzSZd55xoA63Ntfi0yrcwmX5sKsaBGutXlO72L
2F8Kt3O8N77giPKafL1PFUMBhveYTlRq1LQP8B8ZjPtvV05vgE5Ez0ZSFbhY0V/N+vohIflQNSkT
COR6XHf9lDUBH5giR56EUnbKW5sGPCm3sSooinvmPeoLq+d+D0JgQkZlhW9+nHpiEwo4ZiyQBqhc
iy79v4GT8+YY09i1DdkgesTzXuY4IUsrdBoTx3FZKNJcxQicpFk6AdBweWoHodTdfJJdW70xL+GA
ZDEtxifyqcmuubv55CGtCVeKnHVFiyuIpemUQXKYIYuLQASc1g/FlXdNq8M0lQrjz7XB7uWT1LP1
J/Murw3ARhrq+cZhoi4Y1RJeMALNWWg5gSutUFC+tan2jltaOHEkKPrPpxhxU7fcGnRAgigU7kDa
cyScRA9RVC5IHB7UulnIX2Loa1P1TzUPXfuQHDHg6OeNlsuNSvGNROPHKbeanxXv/wWUwBclG+YB
yC4XiCtuV79KrA/duHCevJndtxEcdosCzN5SF0PlWe3nUw+wewRy585fFTWK02Y+s87zR8uEu4nH
soZYSHTBquXcplDPq7IoYNjVoC+nj2D/N4Sz9OIjBPhFn9nKty3XC2whL7ZMqjcRUY5Xvn0uAfIE
skZr1/FtbWVqSkmPvSS++q9GhTOhkik02aNq20ZoDJNqV+mpuUG11ZokbO8KuZ7N7sXkAT7xc+zv
5UKvvNQjgdZ8ci7jjIypFlIe3ft2yCfo/vktXVEm63JfbmlLOHcKNGB6wJfZghxY+BaqStv061BZ
mWlzRE4IMzKkLiiQ1LLpWEU+1iT+KL+oVDawc2Ln37y98TdiK+Lvh6Z0GnOKarDRDNlg0D7HzPMG
JPMS2d2RUjJpeWiDzrPoVwXmI0zP+L4IW5CaaOWZbROGcXiXyvdFrwRG4/iFKXUURuqfFFRDej1F
ree3CNfxZ6oB3M2j97IoYCtUGRqfbS2Gi8Gs/MnoSCfxmWPmsfZVAyzD4ki/DfMq26R30+DFLKPr
maU4i+/Ild7f9rErQbTBcKO1/3hO/ufKEq9bVgXeZtBEfGcw4pliQOzp/Bi+2csj0jSQnWH6/it8
KEAfEUrO1nlAVFzju81RXH7xVQvv4L5WR8R9zl26cmkL8fgGa2B3h4eBflLT1g+/+s0SLrioMGVY
U0m/vdVuQNFwOpd447g/bsXuXb6v2URlTkS29axEal9UZ2EasPIcQUCuGwJmeGgXZhxNDZNRTu0H
V531qcB7hdSgdnel3e/oIDmwyKTW4bVYVN8z9W445vcwpjgHbr6D4ZxRgQqhrkqHI7prP0Ntz0qK
8r+HDimRmqRjMbjDb9LYD7hXREPfr0VMteXd3gYudjEPZRt9trjQ6Jo7zyrKJEDz7gM0C1pvovjW
FHyk/PS+Ei6tejkfhB9c+rtwR4dHgoZbhfTlZ3cDWoaO3yXKoOb86TTB6R2VuvTg8nGcu1/gsRtV
cuIB29eTARoAJ3Vh7KzMzNGOdg6k24+0ObTbIxn+fiWNdhjd9OJ/IuL8MH/yDp2tnbaH/Y3w96cp
HScKVKA8hDpqwQCPqAyVBTH+PfrcBvkIAq2REEqYSBB1+dmhvi/aDVM2Om7D6aCswCRM+4N9sBMN
WkNhhvRgeuuRN+iUNfpjVMXLZaU0mvVJt1tBsbrg1ns6vl6xA6oLmba6Z5AJ1o7EWAWz0niFlHjb
kdx7bH3sHuz7VMZewHcDlUyWBqfIdAcxCAgCRqq4rYmzqpet0MG9wFNAmj6BYsvvE5iuWCGRra5g
xMG4jmZXtAKGdFsn5SpX9UwIY7Yem7qBZd9WLgRfgQqkydpyfcPG42eIMub0zXICp2GTDmdBW85A
k4PNAtxAX2udO7T1thVAzHXM5mLykgCSe/IKfPgeZbmLvkHdYiYgwbn2kzr7xPy6t8wHYKr5Ww+B
cwgSrNofAgTDIL5KGMeAy+HVMn7Q2dO1JP1TERAx6Zr4LhERPLTdwlaOrfCgWFzWFxkP6lQFirqx
1GkCzLDSBA8/kD41gBqlUTTPyI3XdL4Nxr8+5BbOGq1OEUcns41fHcZKDlkWBaqJ6YS4b83x6/l1
Iyd1e7GrrvSKOJaazu38MkT/yvDTSJ/ybvtKH+W6ljFGmyz7ESllxSZXCU8eDpFenXwMxLB6i5/V
8ij2xO5phDa3EH0yIzbmIgnA9S4GsR7DR9ZSF2bIDO7IMylGCyHWsXzYX/KIV8DChJavzhOuIjqG
Ga9WUlxGpsksEN+XkW+4V2Apqzch4svJ2S/QDqOcJ2V7DYynWlY3+opLjT6xD2QNTKs0dCdTAVGJ
BuWkTfI9PioyemKVQoc3DJxcuDqv3Z8A16dDuPE3AoYIlR63tkk1vdgnDZUPoB0+un5tfUc3bNzh
BkwBFeKRYTHBBREykF1JOMGlmDCASJdxW9UxGpHbYVxF4eR2TNBlQ7xhsRuumME23blN9mLR3lwh
Ea2xPnbf6f1HvYwm0MLMOBUTNpcNX8mZHdrLYW2fn5F+fKSCIXn/90hXGNDpEY9RJqa8GGbgooL8
JcdohtDgsrUG2+zGkX38O7rOJAvZ7IgBL9wQ8EAorwCnL8qvM6k2bcVmTajFs+k1vK8bX72Aw6Ox
xUx5rGyCEN+SjLtENWy/DoEXj6DJ+iwXm8Fmkk/6wkfAltOj0xHnFvlgcvCpy3QRJNK0eEsBypNF
nWNI3tQ1GU4LL80LaG+aLCLor9Wm/gGGbcWg4SG+3kHufGTdQKqpFV5JjgxfLRs8gpjkhMs+BaNO
6tNFToWGMuzWLLezo31pM/e/Fe1T7Cdacnker03STFCFyFOLj5wmL2b+WU7p+Cn+f1Luvo8nfGf4
TsyA5wRBGx2+RJSIdICZzD9I9SNG4fpn9rB0eARwjcYii343tVlK9LOvFhK3bnS4QWB+cgeq33Ve
nyxrGFmb46kXhAJubkz3rfHf6jqc5YzrhPe/ySamTPA5UT2ZodQ62PhoLb0NBP2KAn6MHFpsFPxH
ntB1B5DsPwEv3o9uAxr14lgYQ8VgzLH44rBjmaNoM/YrFtynFbOPBaEXEVSw0Ba4bs3sCRJBzH0K
ZvOErGWQCuk1oOTzNmRlqf3+4nbGLUUHPKoiPq/Ilujj2qko9nJ+xUGsQnBr+uvQdzZLxL2lv2iT
+8jhiM+wB3FkjG9Tza9njlwDikC6TdlTx+0HqLPOXocvvB5O4LPm2IWDS5FyiLkHuYS3pF5F0wK+
/+lBbBjEaajt74ePVlNKfEiRpFM63mEAjyoS+AN1CAkiGaOix2e2zLS2Rbakd5mdSwzvaqNGREgo
pZDxKhPgGFSLukKWm738eJv1jw+A3Y7GL5/2dprHbcdkR9D16z5PUiCaNQktw7lgw6DoI2Zfm1V9
tuAh36HGcpuJQXdM9lEp33Xg0RRYtimo7VTES2hF7yzorkjQrhWvcZLYPArc0FHgtCjC1Cnlhnbw
iIa4diVl0Q7TRu6AbQjtxoWf47w3QQ1mIHAgJSJ89+TS7x2dl1XTi+bzNEZlkYA/2IrAqqYNi5Wl
SndATbfPsK0I9uIiBAkaHIDXm0Rcud4LaIsIqktK5gyO+hSad2mNAiBf4YLpAKNyhVsMrnaP1NCy
cfdQbnNzo7zba992ZgL6V5Kr5LWhSgLSjqw94IXU4GO1KzMmbtUs8tyr6gJP7tlyQ8lVYwP2LTvc
Y/fvoPEvzk4QFpdiVaY8EmlxRv98OLqm7EPmDu1EQXwYA9lq4cHWB+Nrz7iLhVVQh2XQY6plFRLt
9/rs/n7UhQUZx3cCeWUcowtjk5IesqejhIH/fJgrp4Wh2MF5B+CgzK44wXVT50tuer/ACRkdKKf7
WH7ufwzCghhk1tdWm7M41PeDrFNk1bEDBRq+H9xYwpsFNDhliWxSLjjvBG1yyQEgJJopOaF/8FNZ
9zdSDwSL5OeUWGOazsnaebfjngVaKQB3Efw0EMbf0FlMQ1x/tS2UULwWsFaT/fOKhdMTVLshqofp
q+idhP7qKR8+cDOsZhGRyF9ETojRJl6vlZzaHKlo2HCBlZawUK8cGnRBpUWuIdIUDZQlM0z+hjTj
ucmLdU4uvVAPDGPDFaYVzHsMKlapg36CYzJcWFvL4g4KO2qtmlOJPR2gxMcIw37R0jh8En2R6pwx
1jVXKQLcGqe6pvQLMXq9spGoIf7pMz1H15XouBnm7szK2/kU9SWdjWQsOis3AAF5/VSoRCLi63eJ
/i1Q5wbKCNXECkP92DnqlILVySSpL7JaI/4r4gletlSme2bOkl9VgUdgFLhqBg+3eAHxKUZt1S1y
e1lRfqDu/OxB2EGTE+WDAz/w1wNbjGMRUiANuoWsHHQV8t0v5GsOPDiDWQ1OR7BxAj95mdO6Z4B3
0uFIN1MZUvAn2JExRkFPo4AwT0zfL3RlGmLsukwI6bQZSrgEev3h7L4TC1tWl40XS/1I6gVqugtw
OezpvWF86YQK+3lfb0B2tQEVASxeXSpqmEU6vx+0BDqAkUoYpNAu+LEzggmB/Fgoq5hJufY3BFhh
HIA3pL+BW14378hM4Q88nxSenx776Ppaw+pi2y4PWM4b47yKZv92WMqN/rxx0bZ+elG+6CisJLrZ
ZlcdVRJsgJnrHuliVKY4iPIoOpF6T7YdlB57HjOsRg5eZAczDnxilaR+pFYYH4RzrLFz0goeiFyc
gtBzbflAD1i4IuX0zanxW0FzSf9kKGx+KZhfjJy/Gz/7JHtX3NsE2xQiLogFEL69kQk5niu5tqWz
LOy66TcC3HYeI3helgR+B4AwwmJ2oLe0g2ANdZNY8x8bg4mAdtFi5D/N3zSpZXWZzIjgKvfqkaZ0
x/1q55yb+cuZ+o5us33fRpcZ2J8czb3T4aZ9WgAm050cTdRcAX5KIOpRfcAzqixtW4Ra+AFChw6+
3DygvNJtsy6gMv61tLsKwAbZetYGyon5PWmXmLgvtA1NUMd3uJT+DF725oouc3cfR6F9U0RYkosf
tYmxbFeKAsTD8UfvqB3WnU0GzEJxw8H6MWdcWBv8W3Gv63M8DQ1t83qxXJQfNb2sy7O2g5Lv+Xnh
+KxL/f8pYj4aVQ1bxJ1E+2nuh+TotHKb78ypPY288XUCdyBxmlt1f1bzIvB/XIwEd0V7mjQi1YGm
pg4qPPULESTywuVfFelWcW8JtfXVLgpsHKLeg3qJCUlQjo7Ol43RSJWD5drgCAc/XFdhuyB1zC7O
G3jxEMRlcICvB4fQweFH7z+gZ7kAymYENrfEWk35bTrkf6ZSrHhXm/7k3e09GoEbl661fHOThUrq
NIvGflL405YtsQObaiHWFEVJXu/mcryTGSX+YABd19v5BDhEyFqlCqzCFrPKOL9sLHbHdnsFFldd
WyJo9PhOpY8Qs6+VzA87SeFfmNfP02MMDyX6cxTJSvWZ66RfFk0/l9BFBdvwSHRHdEXfpDrrk09c
WENUvH9VBeeZbpQ+bFxEIkmhbUCdOa5M6fZ8CBZy8qqD22nj8hJp3j7aedJS38si5KXgXXYmW08w
31A1Tek1+utFWSbIvOiyo41PzfRJZM7yeX14Qk62cHsgqQkjGjJ6ZhbiAnZzeo8v/GDBThsVlOzr
DGhQ7k803gsLRn2xFUC03jazhdAnAHbc3t29aLzjAoAI7PYtnDF3P07kiqLep6NHIMvPDFmEuE1f
rfDZR2F/5Byg9NAXD4VGT6pth8FHN7V8GhWddln6Rz9ir2JbI2OoPxHMtIcsExSK7BlJa2Y+GXdu
cJtAzXF1hf9el2Ikxd4EHNz6n6a+j1/p99SxG4bFuyJHB2fFTG6oRVQH+3o4Vj4mpQpe4M4S2tlD
/oivYnv1y2TZSiep39nWQHTRYQAuk5fMnp1pe1R4oL/95ZZlr6HD9sMpTsdoXkYL1kU6BecCLJgc
pgdNleAeoI/lDxrRfvmAC2MfRDaJSLoNd9Rl2I8eNfAcv3Gw4jxdA6uEIIobeeiwk8OK5RhraLMj
ggpbwcqAobicnHZA9JEDylVOZ4pfs2uz5mY79lREx3qhDXlcLPZ6jaRIik2sY4oPdpHfgqXuWiwf
gi+dig+Xh2CG9U69GMDRtKNe89iAm3H6Tm/qNrO0Jl6U+BeF8X13XRSFKFxcDa7TfhL/6Bms+uYB
GciMJ3eWNcPl3B3Uktl6XGI32QPfX8eqVGVfDj6B7HnAF69wh3YrD3sTxti6ulTrUL6x2UI3G3iP
GrWTP2Ac1BFhnKsXWJeext1BHTCuPALAQzWT8dgcEYPWKYfl2tv2yFl2W12ORd98xVIOyNHgSsuT
9ZsmZfxoYZ8yPx/kWbzpj9Vm9QgTFq9gOcDLFFDdLuFvihLoDCglkHL3quhv3ZiTQILbi+MOc0Gw
b7LPWIy1e50MCctnQQsAQ0EguVfBlgOhRx3w5jgsoJms6X65Jcx+wLQaV846vqkWsCMg6PECn/zg
qvyWSjpH0Of+8ilz0b2yjaCZPQH6XHGTeu5/dUgPVBln7uYs7gD6zxzEMypZc6Z43q5Ot4gx2NOV
vArKMKhdLPMDgLgWyfYpw1SPC0+HRvnLrAY00GOSjjCVzptxYzyqbZkF9If4HxEp96w62XLVqL8w
gHEHkuK+9mPlYNvjD8xHHPAjF+MZheSKZbVOeObMnoJcS+eQ2hUX5JJEER7OvMwmMG2k13Z9Ax/B
XFl77fU6yDXQ/2UGp1a9hevbF5qDycvF4w0cIaV4uvi+i1Up95mxaD8Hxdiy0TMeL3ZBF1j0xVQX
kzhVAacOcx2efu/Uh6E+KVFR7zMnRtwDB+L/bwuft/1XFAlJQMOamSsaxOOJ95iFU2kqAt9LYpgT
tOn9uVGz0edQ0c9kMa84yVq0TBoSg53StG0gNkuoBt4N55p3lrHuUpffVmqJ/38Oqj4bYLMaF5s2
PrfZU8lnNMsTq4euE/giCbxKGrWC2yX2VBoiejnzYkNizjt1AcqvRj45Fn2hidwCIF52qM0CLw7x
cPAZR6jxV4h5T1MJhq1n7J0GAbiRIc0/hqXUjIyesxrJffIberLhLpE9w28FgXXthmDJGzMETtsV
ASa/e3g9lF/Y4DdLBdigHhPowUka7jZ3JbK4gmsM8kzOjtPQIrO2hqvvCprsxL7sb1iSyP52NcAb
TXav6wAfgR8U1D19sY0CWy6j16PNzumGhNuscqtnHhaSEuC2DWBMGFFmQYbif6HG7Aknx2Kdh7SZ
8++iKDT0F2rjI/3R96dGQ2hYZxATtXMx/SJf43293IoPZT2qjNGkKDS/tnsMKvu7oNVvumza0FX5
MqE/Cl61Tp+le06d6z0XIWdokGsChqO900gb3IneKJsW7MQgbmwAt9MyWBSzn3IC3z6n2NgHGLPT
lWU7ENQQH3Cjj48eYbiIwRMvGNKSUdMn33iiJoILthd6d8MjORwDsVbAl88pdSejNI/+i3ufDZg9
wxOgr8k3lyuYz2IKEB4TtNzj6tQMgnZpySoNURqMJz8/40S+ivfk5Np8kXUHFtnYCQ986jmLxiLQ
QNfZCA9vVCJwOqxx0Gr+K+moDqKB+RG4FhhqEKFVZsAek7agNO+9mjNFB2YOIJm9iAOEOEeVH6o2
cgIl6deS1lU4Vb51gQ20mTrVS8yr3Fg4ueFSnT1FvCcdGy4emj0dgFr69Cm7DY7DFIqvJh+jqytW
sCcUDPXXNrtEy1ZG72bA884Fk7cfGAHkRFBvAGMXeZtZhIe2L7DaI9MYKYwCcBuosm2r6HhSGisI
AQlhKmXxRDI/oae66WuJAYJ9k/3OWzHjlBNnXyfHbHWY8bumzE2wSSfo7BsdIP9fwH2f/OqCVeyc
eETSj+wseKa9ouJ5Au4AmXnAlNv0numZQlw1xKRONG4Wj13qWXP1y03GRA5Hw2EYjeHzZ0LuYluU
GNxj/0GAfuB/ZYIRhxyOvms5E5BejLSzkPEaHKMIn9XGhwHYrR0YIHRc4m6+Y9bYLRiAUjvCOyMo
lUk9HnmQqm/AuS6uoGS4EIcwqLUgMzo064BhaGm2pBzpXbdtaz4kZk4dVG3V0rKDrkDuTYw3iMLk
VYk1uc/lAz+BBLiflUAB9HzMU2l0q1HJwFb+IGVzKzKN0bFLHcpAGv0Uz/0cch0+jK6uHW8UkrnS
uGrjtveSe1bao/ycvhvtUZJ1hvSlIwBynnKkyCXl6QauUxd3iVKW/3rH0av+yoHZuEbZeshlzDXT
iBoek6wUj8pt4yexkpygg5pJQs8i3Xz9h4hXntZKJ0NODuNIOc07zo7g58WAsZb+8PVa9qfoNcn2
/AlpRZqvYBOUNvOdwhrvk5dsVOEJj60sn4+w2IRpMDJqa7czmqwMuJI2Igt3h0j19wH3jmCuZH98
MzUB3MoqrbZ+pp0nUixH2E7ViWmlAmrTlhOC2v1h2VtlBSGNUFgd8ekARPdsicFJpn2jyij1V4OD
d0bbkMg/Pg4hSugpv11SAufRR11jXGpZN1htUdyZPynejjlsUjeT2T1UfONCc31TqIyvUp8fMnMS
iLMBcxDVsoSwpACEpALmvhNpRZRYNOWDtrpyh6N2tkwRN34MpYdqFK/xXL1ZtUuXlJSYtB7mN87Y
yI4UbPovc0uoVoU8lk7mU1FWr3nhB9u2sjLUCKixlFD8du9g3+KFg3HJrGH7OH9Ah19nTd+xCr+P
UXTOqeBdICckydoTZrNPGX9brtlpfiE0Jq2c1cue5cbDXtNE8s8oZaffHbaCHrZ0fvnYNe5kdvMC
QoFHaLOzllP+1IJt5YVjz0kQ4HdYPVsnfWWwlQmDvYgnsvqrTzmoATckOeqdtXmdZu3HIOYn9oaU
GY5ZqiDt1Tw7dFymRl9Nb2+9Y1zeTKkg58z4EAfBfXw8K9WRGQX6oHmKPiA1A1RVaOtE4j5ZOqIX
h+MWjo5c1I7T+cyWYenGGGYZ06C4/M9v173LQJCR5JU4vteCxa3Ytd0gwvE97KhyhB1cMAKG5nV6
jUe5PYfswafpKopUIWZ/GyRF7cwQp6Qmg3ejodHExj60W/wGMsN0KBsspD32AcFha+2cJrx/+90f
ZOjAoyO4CH9F6r+LjC8Y6mB97qkTCrm8UAAl4G4xyA6bhg594D3bA7hidVIUHPmryUla2v62lQVq
So1gJFKQiilZabSaeAfNfXKpwd2SoMDHxnoIOqvhjuovoZBcFb//5VbMKCB4cZ5rsjAVQR0ZH5eB
fAd9yKkc0CVh1DJ9GC6rpG9gyWlAVKcgA7mBKCsEemNn7rnY4wItGrRF1KnLF+6fmkjwJGM9V1h7
qlYsCbL1s+tYHos5LfzBEwl1A4pFRWEjdxKXXr/G53BRdMjwXELrsP8atIgxalesdPl7SdDTCUsE
ZrZE8DHPukzeqngVXeFp2VM0/lLH6Qj8KmvEsDmHhfdLjuh5Ak5220hfhhkBD28qt1DSXuh5U/o2
fGNOMX3wnVetM6iYcXUDdfXiyAcrxl6KgKzaXDwla/gx+nlwbTkUb1KJnruVvNh1jUpN+WHGT2o6
jSamVVbFhUe8J1VtBAluiURWMWSbJW7CH2Uhnh6YoDgSQCBfpPop349Ts3XBm6FHFGtEN+wZyL0L
hibTPx3YXKpnQTDJX1kbq0Sf/6TLSoIHU/KP3lyS5iuVAdzKyjnsYgvMDR0qKFf8yfVurpYM6/X7
MOthki9H9B1y8gOVOMxfO6xSZ//xZUOB9mVlB6ZUbm0oi0Yyp5p5EVxE1iMDD9jbx/c62GbnHt4l
mrPv4Jh/JXkA26pvzUrbCDH1r94FZmupnOYFOaCfinuSg/BMCld5ZzuPY3XDoT3vuJGQVXEp+boQ
rgW0kGvmAznCUXjP//Bi1eWrk9fvOw1L8Ks0rM+PXeOQh+Yu1YZvBgRvgUcw6t67j+yR5lfWYEdi
aA2erhvkUKL24uJyczRIWGvoMSBrITzGVmDITgmdjjc65Dl1gQ3/KdzcDArrOKrbQFsblX0+1Pot
e/SSnLtjAR3/CtxxSUK2FysWHhQXbU0DAQqXCTq74DLbOcq5Nae/P6Q6bPUGBSTYFh9vZWwNXEjA
D/eBB+9wI9kXdpKT77mqzIGtHxe9/S2YT96oFIGDDThVrlIIf3i4uj8IeQtuiBRQFxEkyMC/Yi9k
iMvWzC7qaCDeaxx69uYL6weU+JOky+ttRsvHzU6XGgYgF7kdRFmpJkak2KWtqCdbznWUUUuufO3F
IeGOQqfU1nB+AwaeUeZdqEL7RTLCy3ig8fv7GSUc+7xPAJk0pYBH+YzAGFhODFxPBJJyS6RAq928
0bqUe1p1/kuTQQUjjNTOfyi0dEiZH2TlzORX31doXfnlbJQK3ome4HWj+uVWs+4dtpYevXkuUN+m
aKQtngPHS0svQ20nd/whwg/CfI/hCvDmaJ5OXJj8WWN4bM2e7zSb41gXjeTkefkWMceDyr88vg7H
owjCsJ0EhTpcxInjim9CWW3X0dEI5awNCCGFLFVLTpm8+mZ5BNOSv0Y33vDyHIihn+FcuOEvbBQw
ce/EyYfRY+1J3eAhwUm6NDNXTgOF292a5M8sBXq5+/q8PuQdBm8H1eB8mkOWYtcnIltYtXk5WsV5
9Pb3zMzQmfH4frgau7r98kkEDUfklK0oN9Ije13ugCRhXG8LF5VKbnVHVkJds+pjrZbDwsrmpAeF
HI3nz1d9ymVpIRLmcFhun3R7urcttVNwtZLNADnA+JrAniopeCq908WQVuexnEAbDI04M7+l6vyQ
Vpxi42cEioWZXKSbTDu5OL0PpmBhkuzzrNjVCZsPxff5TcZjviPv+4IB2q5cjOaa4/IO+YzkyLiF
V90sccH4rflXF7N0AaVJfdkVKIZk2WQYdxIvAkuu8cG/qvH9cNfuYIOt6glSfFLHrO91mH8UOSyv
DzhQp0kN0n387UzsPV/ffj8Ef9ajW/JJAr8sC/T7JNAHcpvwcwk+p096LOfv0EKhomJOF+r2D8Zi
Hejz/FDAbbQ5jkuBDRsocL444q6fVUoLtlM3c8AJl+tR2Zwm+c+XGOFWcloSTNL4yPO7+V4o/Y6i
AI5GDxxYVfcNcFimcN0d1ZmRnhy9nP8x+zjqd3RdgLpylN8GUB/laAtaY2ARgTKnzeAHr2s3WYK9
rGp2w7J4nIkV62uvzSkmvf5HaRIanLkKB6SyZ+Lapu8xXbqcN6s0xOzCgnGZd7jq6Ys9RfJxVKJx
OuSmDABFxEjGbLpEl7cCFcK70IU9HxCvQnOofeyEh5gN9HxUDgKRHfe3DcFJII7fqa3tTK4ePh0r
ZHrRPmDJJWfVwaY0l+zLO4u6NWp0p9tH5ljRsgYAT7YPTu9QTVsoLaepIIfMhFFQkYIJMgeTQb82
27EIbXtTubguhrBgsuTDMBUez9JCfyjKd1Rb968UN0yIji2YUlKJBhkAMIC2rrPXg9QulfQDkhPK
34BVOXTv6DrlhWtc6v0m7SNSQko85IvTi98cWL6lzN1z2YEwa4chH4J7BRvTX3sHtCQp5tBnn2tw
/DJkUc/ZP2GqjSwi/4/wp1xuqqWGLtRjW1rM2dZRvlR6qbvS1LC5UsJ5wwibEkRItQfdWf0nbpyJ
hYKWASRDMlpfcYIhGs4Zwe8F1fx66aaCcL+c5FHikgxLQVXvp2GgdVPjwLLUH9+FMfPmO1KIbr7y
JedC4XfHTjC90uOxKlgZuY+YIdgd4ob830soDIlYeDzOnMVrMDMG08Li58cfMq32cK5Jgzk8K0QR
AdxIV85TQHOr84nHGjmwIRdS8xOp+izLAF7/39QYXUh91vPjDlp6EanJndqeKSO6S5hnN30nT9jG
A3OrmOqFsl9TUmIrvE2TUXjXJv87z5qUogcW+nEGJZYW8IGZ+5Wobk9l6VhXHgWGRw6PeKF3kJvs
fQDtf4O7MeVRAbV1PjGQKH1a8f4WC+wgIizwOBLFzhd1TbTZN5tTfHmz48d3Za4megcgX0Io/L0x
TMBDLl0fCExXk3WY15MU/fuMvVrb0f96XTO0anonbuJ7RTgtlIi6+nvch6oeaO2C1lZ7wqjMFHNR
3ESsuYrH2pmTGQb59ZYZfMuSV2vsQT2RVXyUl0amZwujACKukx0x8arau3cMQNux67jpOlvPLHzk
+z4MOj0N+eeN5LkHjrBFoNvyd2kP1e8dalnfZ6lVr0nWOA2c8kwnIiemMDdtOMYupJfBkSiiflT6
VkR6R3WRpRp8R8bQq6IVe3c6qvQ2eyDgChSWxmFJseG1a5pxDdkuauTkO9X0YyO09b9/T9mk1AXW
qJRKWV7Zq2K7ASOGB06l0GeeY5x5EIBCWhy0iFp0sV8prebcYzEMn6glETt6Qq1SmSI4fUCbBpre
e4nWj0uDP4AN6XVBdRjSWdy0D0jIIhS2GIQu7Nsf6Q4bq87gqI4ioClneSm9m3QZZF+jGUupGj+Y
HvIHpEkXaKcccewXdgpPIWsrLWfZXUBXWQkK8QqM6Hj/vpEjD6LY09QwYwmecPzTsOcppXHRgIgq
L19xvatoUl4gJQe5WJyQ1K1LHIZLFPgLKnO+D+9GRnSIOJRjFy2RlyIVSEgKHyr1bS3rEKRNNK0a
Glzthie5798uuJ3L82oRV1PbBtV8LFdYgIlTCCVghd0zUirLaNWVUey7yoOsk0KxGLWSFyG7mOh3
vb3lqfJUGQb8FSzt2Rhhl8aA764skj42eSu6RoGic4yb6JfXR3JmxzFisyGya+FCbmEc8p7sP7ux
lRxoNbjMgqC33w/b6bMfv2SuizBuwrKjDH43SuCz/aqc3WUIGOD+KKAbgv9Zc9fpAjk4Vb5/+yx0
933BtbZpLDWsyhjDzzMk9q8PgtOPLRC2qCu5RbVN0Mh87cK/K+J4H5ImGqrTOixLr8PqSuRogfYs
eJpZcQenbWZ2xc32nIj5ICdgRnJGruPMiCySzQdWtT27+KBu/SondTnelqxuIt7o3Qdey4PsSZbY
7v7yDZIxTBd/IUvF2b7W07khfl0SrJlg0kJH9WG3LxCkNDdA7DYKfgXMEft7PwseYRprkG3KJZZh
lfLvaF1XCO0btUW/OrY3JINdTwAUHaxr/XkHvaAEkojc9Umf/tuiiZ97v9gG4QD0ZhhVLpczrsbw
EN21wcKxGd0jnRr0mK10iDhPkZva8NQAKXCwdTKijK02J3fT+NnQSOwfCKPFqPH0yacfNfzRQiXs
uEqraArYdPc5XJmWmVnnBqsHQJudYEztgeFnGimr874YwfF1X+YILo2CPTacaEXpfpXhBxw2XOhX
NE+lqVZwl7yaaYcSB4c6YGBoIThGjxItRRnyCRZbkq4rF+tCvb4rkqBwuQ4XXFOZ3+gkfIDXO/3W
oC1TbF7OIFfOiBJiiWsCi2yfYGvjvOMQJm8c81gmKmHnnsVkJg1QFjDtszGwsGhHe7OIVnsdPiwQ
vaaTKvyT4fimp2tX2N9dXHxktVekPY7tRv+PfkUHE9t+fv+B0cQJ71GTUBsq1B9R9k0+1ePsicNg
E2LOrrVGEtA8+SZ5zauXLT21msh8u8SkPb4SHq15lRXzeP9cD54K/iLV/8GmjVMOiuFD+4Lx1IFq
9AeO11yr8/4OUEHTDbkPipH8P9q9x9vPoRzZpmU+0BfbizaT6Zen8ZX9YpmdIPrptEeQVKDC6eAC
80cGnA5jA4zkG4WPzB/6tYG3KnRUpNAblWVZ6udeqkob0AYjzA+W0FN1YlAVKiboHS/HGpMlkiUn
RAHmR4IUH8hIdHUV/n28ygx4CyzCcOUxNDIsGJlJPBlvoYsKAIIh5iBkKV5G2a59I2e6KL6LKPrS
Yo20UJjvuJuDxYINXl4gyW18HNiFXhhw/3R+5oD/vwvMwbsjCdQks1stf1XNC3/qqhbexGDDRRFk
u6J3kidkv//bm+Z2HTEeipjvgp2kB/MoF8CE8XleGFgIlR4H5w/LOgHEqKneXXNx5ex1x3itDhvK
i2HHUmi1mGG5wiuFvEOkEv94oBjlNx8MR8YEPyMiJSnFoJQsYrVZ37EeNN5IU93ZULYZYWKShlyc
4nOY6vJEiSN94VPRUPdPMZ3UwzDVXfUhC1GHp9ioi6XqRtFaPkqiSu5kJ5Qdw4gRUNG+twi7OFko
aEWrk3yCcOZFJFrjKviRPP7nt324W5pn3KcXopVOIld89FOPtSIxzryk3Bmk2tNSvLTIqtSBuo7u
esl4ywMlYHscbgjzC4F+LAJNB4yOmT+4djwqUVfjKjQYGhrDbGfsXmnjleXsLdG8dAktCxrafQAd
AK3bORdMNsZ+QJUT3EUJjZZ8Pyy7lbiND+FzMjg1B4bHkF6XLYZ1XZ1xT49B7J7l8RxH5NZgvroZ
zIhzlk1MdUrjj8CKqPgiuMhqFnjTKS0CfXmabhnW/PQ/AcaZl81RdDzwZcFcrRU2OatK2XSrLNNz
CubQ0/T0mWpobJ0DOWiK1ZJPk91wZw2WK8tNnHLPtybR2hW1b+CVyZl8/rLP6DeRA9eetD3ejEn3
IXkxHIMdO3BRuz1Z0lAXciJcuWW3cNYpnmuRcPh+QnBp70oAuWR46aQe5FSw/nW8YyYOQH6KOnsD
ohKMA+SQ5CDjspJKkmhknRkRRAxHPJa+uNw8cJy49NF6fZ5tL37idG/rpYdKpW2bxHxgIMnHIdFb
b11r2A5y0YSCAcbpNqC4eV2K9Iir40sglYrh112oa8h5pRuSIwC9XqCiVaHy3HnO9WFldxSSzuTp
82cV5AGc+QITe1zjmAh+AZtB/GtX3IHS+4t7lvGBgvHMzYEnUkqaVaKJk0ds1zX807Oxey1Wsekc
PUeD6eMyDpsEwXVfoaS5g+IKr0Etr86dlrqz3EVnYeI+wHpYWhiLAzFovwaAHUXB0xU4ItmvX2c0
7ds9/NIbxy5Pb4SEZLyEYp3bTcuGcvjmZLWMP0/tZDvQlhUHtT9TBrWimaIheLMC5O/9CPl4jXa3
bdNy6vjz5b/zZl0Qc7binmuU43517d/veQNCX4iM16d9B7ygxKOP3DSppyut78BOPjC8g4p+4u4S
chrt1tS0CwBLLsm3n9OeHh0UQD/Y+QjJqhxfa3qAHb0Iueqz0iRUnDzlEbJYN1euhJOROv7R9/uh
pKY0ThfV2mnrb0/VufQ07Dc+R5RG9KC+z5h9eBTeBBV4Zo2qxlaTx3XlqniZR2GOimrNxsVAmuHl
H7nWUoeN9dTB81NK3RMqBeqB1rAbLRNuu7IMfhDbAHQW8F/uvsRdzaQENTdVheeeevVyYHJsCoqS
Qbw+U75/ztImXzvVxYm6aK0Xe0IHORrNVq0DrUcjDs/jqYq0NWiayn84OH/y0XDZ/gIAtd7WQxAd
/9e9sIS4ErKUrUfFNjEP6SRZyvDpv27I8xSlekvi6MfP4IhuzgZPLDX6JNZhiM3WnZifhM7IauAK
1A0WmklR6dtHrFoAaupZer0AV7I47IozfX2tL+ooB5RLs80bjjiaCFBxCPC3HHwUNRchdT6gEdhB
hzpMb2QY6D5PIeJlGP6U0YN7g5qjowBGa/K6o/yZzoEQGWtw1gauONvQ7D18O98W1J8jfRqW5TRq
UCoENPqvwKVzxtaVsEdKQi2xy0z61NYZwBa9x92o5B0rpNnQ2GKgWlXC50NOFYjymgrnJ+CuyRrJ
DK/aX98UxuvC+JvRMyaBtGjzkjs9qobbcOSH3VXSkLMkyop8Qn0j1hOkehp3V73+w9/excz5Sp0L
u7L2LkYSvc9PgUIddDO/QZU0cCSY1B0qCYoHaxYF0zoqZN4BV1t6b+wDju0cm9ZyRHkHmpu95Xfv
3ouOPo957fGmLzVtb2Sssenof0VPqxTepeBxLV01x7rwnAlf9+emDZ/xqbOt4ozF97dOCAKjfOxG
rFavy9DoJexGvIPz2QNAQ9pb/M5t71hw6+go91GrfkUNDYFtoE5cmL8P3cW7eUijGrxyY8R3KNIS
eaFTmYv7MVn2uNr/ueKoiSNR4ZeflevjoUFbG+1Ke0Jga1TET3oKUaBRXrVfFgN9sKy9qnQvcYXU
Ci9hkFWxMxucyQFoEqZDVGqgmpB/y9p6kCQV9/Umt+9dwqlvtwm/7W3jnmleIzXpJqk+58O46I0g
A92gAmLb2riF0Lk+nrO7Ny3HxmsQncI0EB+QQPT8E4hqyNNnuaD+RGwPwXDd4l7kd5rDdqsnFoMr
85PSlLxNE4pROrVXVTmlVpHOZ4GGad6j77l4k3VJ9O6YTcpYvJjOAfZX5Joz4B11+g6FjNQvIpXv
sJucQS8hGK+Q9E9UbSZ/IbUyXPd6xTTA8FgWqz7YkvCup6INV/y1Ak3pG7UOc/xtMFnFAOHdlV2V
jKIA7Uj9fE6ped0UldupGNSDQ07r1V8tclg+FVhCABgtRmQ2KUNZrmkgZh2HX+rfi7YxxQtT9D3L
+K5NR+fFx0oiHCWMjpOqXVMmcx8uyRyk+yorK1VrJz5wGhw9q/Yc7PH6PMWfOBFPzk0ZpgehNoXb
PxWlTgZsa8uM612vKzBfSOKaceVFFaGWIJ7lpNnBm+2tgna99B9BTXkmUKKp5SJWoSAiteU81E4S
YoAeho6Iasx9DFF8rEiIRKw8khmppMWa+iyuv1uEVvuuuy+bbJW2Cwc54CC+GFiAmAgBtvkgNTvo
TiTMyZWPMDdy5MtND+2A6k7FRraMEXOj4Qq7LasynJ6LxhvWQRm/1uQtQQvtro/5ZdzXQ/1Ow/FS
BgI/d6Qpeqvpmy6V+XIXk63SCCQEj5TN1tZqMyrGMm9XTgDjZt1Wq5DjzB8xOZMah2d/hbPv2tF2
FVTrgc/K0mCpttTdDIxiYmgMuodOgNq8A5/0syX7P2El0MyUkcVSR1kqtYYZ5yuKdllrvcMxgBMJ
41vwJqDWFv45oJ9e0Wt7C17DQpMKVasZp6rdXgljVqdapYYb3LGtAC9rxUZ7kzG1tkLOjvxax+Fy
OKnfqvwHn+fND7aFX2B6Xnozi4RBTgmn73iUMYTh2c1jhgJ6EetrImU9dxNLB3AqoA+IiADLYW3W
bUavTQzbElfY4pM4+Y9cPQV5MnoBSLqcZdMWB5OdggWLq1fKTr9YvACKDAeTq94ODBLbxYdc4nIt
+ZcSCN1hvtX8TlN30lIpczFCabyHdUTp6+ohVbW5jEVxtsInDT8YIkrKYbDGdUFA9fq+PMmm+kbx
GcHqOHPgw6jGWDyhbfDkOH1mznUSqBYurL9bgY6Z14y2GI27IaEeO+ihGkRit51kTGUtUyXLu68c
hD4zilAasAu+2XqBtCfHDFUNM9vwYVIW+rzhWX0/tN/iHD4dwT+35PzKLs1hGCGxX7d9JL5N/oZe
YGnhHYKwyZ+pY9Cy9Q/aJ3dPTXAZCACzIIIBaJxtxAWXHg1DGkBcZ68+iQlsiVXn5jPxfUSf4hC6
LZoJvrbp+FvNA9CsVQikpEb3v0VF82+PHHrLcaFnHahyHDlfX4590u4yomPqGfSFxtUMLSXCNfvy
ruOdYY6EczaQlGMctiibrN00p0Q9ZGdCeIdr+JWvlAIxBAQRZsFhGLnXNWEFIl5MretZKzd9W73H
xqKxugiI2+xwaFPIl/bY5XhuucwNU9+OUOfCFtL8ZiNnjeTsxOaj+5aTLgr1DarZ7X8sPbHA2eli
Fcn2V+/LZO4QZD1/suRZUvDpLkI+IzV7HAcFulj46NqwKyw4ROhF9+jPFU+JNNYAmctACig/h9XH
YQ4EyG4ovNcBlw1SLQKgej1r/ug+uy6eLu+1puOhXVoNAXdF1jW5CAr1raMuZobDy2CzJZvFg26d
QPfGwUjylP2ccY4Hbke+BmRu19jqlncVrasaCG6SZu39+uHpkVBU46zRpeDe9DKc5ywlzRnlTRN+
bF0uDBBno9WoUQL/3XRfhPGDxqxnHNo33yDj49WZp7+jt7AhidYCRrTmH8BUc/yM1oVp++g68mf6
DbCPFaY2aUHZKlZhkeLTV6uh5GGOkB1S7T8XFwAtL94sVwo1QDEkAQ0O/rVxVba080Q5EpRkNnXW
VpwdXMHxx9R0Z6UFcLUkqkDNV0tGRnv5WM21DCwkQeW0FKMvwFdjeiujMpFPGO41eMZyWLwI6YSp
8F1k88MK+7iNCRN+hNkxwLKrYq6zGQtgVFUoCbIBkzrTahNR6HCcKbzFffOzu3Cj/pmXsNaFo/GZ
kSsvCqWQOp2ELGA8LZF8SflOuE0E607OiXzHwczezrcJB+z/xky1pnlLHXRN+5rLDug4Bql4RLQ4
0O3vE/kijoGBU7LqORheHSydngVsMCewHcQHzAvyecFrg/sIxGRm5xRRtLq7cQIjAXMGACztoc37
D06BP0LubMJep4/WT9JG26NBGRB1TquKmrp47ZGE/hcs0ZeuhUcL4u5YUoieiVzqdMi38oU2hSSl
7Xoqc6F4D3iu689t7gpbx21tEJbwFTf3fJ/f26TciPYTM44c0VLnd/xihBjECsOxp03dxgZNLVDo
GVlNCBLpdAS3KAYeO81Sb4Y2Oy7gYkJMv0/hW1tNL6TG1iF2Z88QdUOIKGB8USEjwCq1E+iJQFBV
wxUqRdHFjJYDwjmy2BUkhPyKdiD8l6H+tvSxu5c9VFD+2Hiy3aeYNjvq5oTpvdnMCffY6f6bOdTK
x7NR1JLI6xQjgGuF98668A+EfIJtW/xXu2XbxAku8UnArIyPNcj3Opxm8+aM0EaOVbDe1ktmMwce
T7AhJXfAivZXD78HBxIqGuK8OojAd20wNz7xbmvO8Piy+Y3zAnx55kNH363ECNLdlydV24DSpbSo
8ZtDkOlYwzT86BdBfVdWnUSOSTPdWq59jP6y3RdVoA52O0u58tIzrAy5HZI1mQUSjQH6tFkcFi03
aA2ezIsJy/Ku0tPKnKHRuqdkeuTgKR3B7odGSqjnhcul2azC7jhAJVPl3u04n4ND21dpVK+cz7BN
t57K0clv2m+Sl3WHqlGe9vN0DFG9zETVMzmz0VzEXWg9X8V8cSgbsThvqdHPu6r/rqTXsNfd9+bB
1ENDbJz6R714axUN3G9mLEnaVXh3xa297V90N8HzTtDurm40hpbbL438DRgR4QjsDn9esWma6Jk8
P1OF0A3yWgWhK9wSnCu1ugrW4nje0nveUsZzliAFsQbt1P/nXvKdNgW1bP1zEL2YmPY7k1cDoZqd
OaeNOycc2MozTh0ijWbTxjngcl+X8TSgGIdJIiAZxy7+ztphU/CES5WMp+EuYULIHHp3PYV3cQrR
iz36zpgACTxsY6SFw9HDNobhPX1OzDDjOWnV+/BD0yDXE7e0WCCeHfMCg4l20VP1Jtx5Wf/Nzu83
zbbCACwCm3rqrtPM7zm9c+QRpEgzXZSmuYcwCW0ae//odkdp2NBKa1elQZqDBlqjsq939Xrr7naS
DdanslcAZ/eT+/s7lr/HOcohJcxXyeGKmsUMe1aRVv9RSR6+Mg+hjL3u4uKAi74VLI4P/SnW/5Gb
i0V4wMkOn8sty9E2o47TGlGVsBi0jP43tXUZVQXET/AygaRgbIoXfBWqlXSMO4KqXUn1L/Vr5UHR
T1WkgRmOZnyu/RB4z3YH42kpnSREJcR0SA0hNdBc1SmcvYLWRbZggbGGW42kB11Gv/OQlKgbtr2r
gHOHPcbyx2iddycvX4l4+/bRRIFSpI8c3St2eiisJzcL2C1QPuvsK80czlT6TVpjVxy2pEB+Uu+Q
Wxxl0UJDAHYM3W30OZSsgQVdbnUW+nmdeQZEgebRp6+Jvz+Bm48sQodKTT/hOpLUcxiUuufTGrWG
q/vBIn8ckWoKWFnHiu82q5iXKyXY217n1INnLq431TonLiw81snlr2hCXYq7kxHb3z0rAAa69p/s
O/gvG9lKaU+uNTTlmKqbhvL36g6hWLBBvcROpmxSmC67xpZGGoRReMCZud7BFl9c8JeeMH9Uakfk
IkK3dEQbTGlhyzmomN34VM9koKnc8ckmce1vAV3dAyUbv2PvJUQZh756xO67MQNgsBgrcXpbeNog
VB4UCvLrAYF86HZleGXPfq/6wARYtF+13HEZzctz3Sf5UgVPfNnafO8A98n6iCoCyR2XCD6J0sic
fwNezwW5Ezc0FQYjQ9htgzbbpRm2EdX+fi5HJv8S6Srm9z0q7Au1TvhAX1firBKLBH1oIb0zMo2/
QAswI3oCLgWMPcSFVh6JlQUawoGqdFLgFMm2nGQyyBFa8CqljzA8jM7lRaB4uNRscdEguz/ceXF4
O+Wfb3IAtLV8mHJWaDZr70xTeacUvH6DhuafFN4BInb6fEOZsCHleMgUKpAjzWXe3zQonmBqPgmN
dlVRs/um7XJkNqZu0rhX1ayidOSMftoxCFq2BudWRKsJXjfO4BlQf6BbTh0RCxBx00oU6MRRS6Su
RZg6kPsaF9DMTtEbGETQizPYa0WhNJgTYbp/D0Q+LJxXCrGjNW2Kxu3EyFc9/JNzWNC7XQEiaizT
RtYf1sjnff8LX9al2yvlaoRxKIjop4HsPY1kgXh6U07dLzAWhT5ijoCRkASZnpgPbVtFu0P04Lkz
IT3KsQ3bxXSIZcDoLnWGItqEYosJ6KmLqXRceA+St5a9s+RUBugDV4Av/0IhXrwBt+Kk3cSGK39B
rS5T+Qp6xqQmOesezgZmK4A9Fm21QP/iUfpeR+CwBwjtyk7ecRwz1ZbGjVwyXLOUWIej7DBw68dc
UQ9Nr8ovpgr6UUCQMtGbhlMpefy3ksaCYO2rZhTPYBBsH94WlnU1F37rnvmBRVPcQhMxz+2s9UxH
PguBvbwSpergsfSFL/4ctQbYQbn5eyNL6vJzKShfEt93pOv14axRqD/MlRXiLoC42/Aq+S9FEfTe
ag0D8mVIofMXvHDx7DMXBl8PdOicyxAd0DD7p60Q3yOcv0dfpKWW2qM7iDaXiWnCTr1W2lMlnVpC
g9/1oS4aF1cNYOHnnOPONMc1SU/2WwBIiJNHuvAN141hECPWngGNe2Likpvo+Iudy+xiP6aM5KTc
d4/p4U5sCORTRFbuY8bMnnYof68c3cXg7LU8WtEzgxgUp9Uy9RZuCeYLDOoQ3vvqZtqG2NxedLZY
PRYa4vcTSUqU+5eawuI3HMXty5t9rgPhx6fZB0hsXdmFTe6v333BN0BfxBpLIWk6IbA/bErytTGj
rC/bTEAD9dyzjchfBBB5XNY6wFfjchCtPsc9bZiCWbTfefSRMVPb/CM1FY3bhVooiGsU0mds4cp+
lhSJ6wG9TwflyYVfB7j6WZh/IQWYAmwox9H0DUJfv2QcktxGIXPdtmEMwo0uRyTXku4HpgLxH1r3
GfAJ7klQI27GxfdNj75SmV4IYd3ag1OFzr6pwEQIMk8H8CwrhJ9j2NIIv65RBVXBFpnFLS8Qm+og
jnWtWZAqkpRRHnCiqRVssQGc2tS2/Kll52DM4kwf6CebA6DJ94L5TtWHFmR/vRHWmaVS/rKcuWfW
iB74Eao5kHFJ0E4tFbLZCsPKKbssh8r2cWF/X55S8YRMtdoOrHdWminSMoaxOSl0pactKRymv51S
xVgFmCryXVkaliizyC+OBbh5ahpWqClh+ZJbhht1t+NsRZpFHk3JoaSLAUM5bOvyAt4yCqG2MdLG
Nbj8CHgLUM5Ddjc43GyBCTm2DCoA9doWtGoNFxO2w9Ny9MDVFZJ7K8Re86DG5f8/fNVdWTBjsxbt
X+TjxVNE8vGsgNPP01i6aKjGRBtr8C/hU+blSxa/zSKg1o/gS8k7Y2JdL5IZIV6glPEPfiTRGdmR
J0EDVAIb2jjmhD3gheDZ8WZdWCtB9t6YK+mRXBPS25jMrskxfb6pNh24KgzbljyrTYjkwAH9JME/
QjZjzAOTX/t+RQk915UdfxPFE2Zz+kFWO5w3Vl0+Ml17jlTeLRaGKPtlor4B5yurrpE/hZNDR11I
fZuoScpmKPB/HvjxtJHyzBuyE2shs2XgdmIL92oPghLHWBUOQh+4XAnSA4zoCmff6WqfDbL6cSih
LaAN3MUCSWP3pqxhI6RQmhJ33xP+FW4/XZAmaIX9Gf5H553r+GDC6olMcY7OVfLWl+wOVR5c8cuL
c5fMUwmK3XyBjNwoalUb9lnE65eIX315ob7GISJVf+gaJK9yOFhISfGVwJg/PCCohjS9luJ5+tvA
0LOQExbRgr2ZGakVnEq2q5k8zinyRKCtVWIZJ5ZhWCiATWI7NycnzMzZVYN9vAtZ933AsSC6Fcud
kt3MgrLQon3vVZAlkPERVWGrUxlK/8yt7Qf6xmCYlzmk7xicS6BKAho4Im2O5CV0yVdQje7lj0NJ
sliJz46V6vE50yyNd3r0ys/qUYOzCgEhzvvqi6vhZZGIJgsMafppiFOxIGdpd4CugAZ5D7gN2lgE
BSxv6/yMcJl01AcKB3hPWL7u7ZwFLNi4q/Zai5RxAC2rrlsAZqJZA+WuFcYmK1mjuDNmnLvU8C0g
joeUPtU/b29nwFaVPE0oip0VrJOfNB3OepRKt9Eb+welDPPro2XLnHABIVEbOKms/6pJbNV0W/3g
lsuMtf1y6MLQ25/DVfoObqvHCQGPdR1rQCkclKUJI+XaGHvHvqXZ/df6yWXUPzHLQ5ElLOWjW0Jz
I9R2xhZDgQGL/BrdDlH+rE7dx6Z/4jLMyo8XBR8lJMHcoNIJKAbvvgA/RCcNtd+bAymUsFeaEkeK
pneQLwKuz3qf6nQVgZ4tcrpT2xF+okoQO4KTwMmzBf0vSNqPO9oHY1EF7UlxwcM+dai48H5BTdEZ
y3kZ9KEE6k/ztO3i9Cp/BuZK8nPbP5Ws0MSWnhIzcPFTDl4q3pYot2BbYx+nmjQ9/93VlmU2BY4f
2V9fi1njsPoVO6JaWMW75zGwJf1ilxK7DBjhHcCrj8aUmTxCAiZT5a8YEBs0ZbDhCyOpMyme5SL2
DYiUbiOVEgLY3Q29tbIWS+8O7/SSoJL3X/qPKlZy53cLQ5Wn2iVOEzO23c3GieTe9ENMIYJcC71o
RxUCdXuFMT0G7Hwk5oKDIsnyeS/lNlQ8xXpT1y4iwltUnV4YD4fGg6eIoEDXt6e5TkVS0HhvVkOb
JiBGd+qAhhzzZ+w+yE2tDZG7iJJCTGZpt5PyyP6MrwNvE2mHUw+ybgcVlOaARnXFExHEBvVtTZPc
B+zCd7nNBsOT9l7UDG2sLNJ+3IIYN/alJ+2vXfByWa81lT5RtTj5Yi/OnvUmjLS64z7iK8kXaIkJ
dsodBYp+Hl0jttUDykTD/MDLQiSAOodwwJC2kH3Nrv8SkP6zkgCBo88CPh5bdNy4VDQDOHrN9Yok
vYRcKRYzvGIqnngSiWLqMSUdV2lta4eM0zuEPocc91qpdFn/Kn0QCNZngdl3LuYboGkHZy0AtgIv
KNGjE1+IMSGlTT8poI5Xo/PZqouN2Q8nc90VGFCoXBJLrMbHJAEyw2SSBzOiOEqBndaRxRt5YF4O
5RGNFxgQEh4/vm2M8B86nemc4TugjcTY3MeBDkKcdE4PZtRqbz/qDORUusn2Afe3fFcSKz2r+NHx
ZnjuWp71CvpRQU7P40xgs8i3+BjyTrRuEJUTVUdC6AzyEar25YKJwjCasdYOTnW3uKzO3a+bQkxl
5aMvTB9y8+zok0v5tpFEixV8mgC/lfbNKjXd4DCnTic+4AoJ7bmrrpdiGg46q7iozMfv4kSzb02s
oPgRIowoN++zM+3zzv7z9G1vcDfqUHQaeaVJM1p8g6yAT6IvXY2d/3kA4a1ehQ1E37VckLp66DCV
oDElNvRLySEyAlKTschZcvqnWv+YA7M9g7UhH736JjnESfXBURotxZVKCERSgbUMYZkNbOrG0gtg
fNvn+28reP46BVGOuFkq71b4ZQyOmToaShCHZUJ9TMXPnNkiJvoSt4yE7Dn3JhgLw0LavExT6sdJ
o2aItpQIqgpOHov1nzPWKkn4IeSLY7iteiJOrX6QmtmnKFLR4YDOQGnLl02L5CH14flInAxMM2wu
TXtbIV1wObpI/MWG8N/tXJIbV7G6Sf46RK7YrqUGJsoGdK1Qbbiwo1ckfLFkiQ1or3LoOgINaDHG
Wsn4bwBl9fS2W+mSkdH/ABa+8LX1yHuZqhI8GYWKLhVZaKU1AvQ2HC1hQ/TZPnY842yGpDHg7E44
yjpEd6VrUUT4oqO90fiH9XOrWrjuUKzv63ej/zjaS+AUuVsVhlHvyds2LYwu082kiDsuH7xLXnP/
6Ecqom4Jd/c+sYqxL+6iTcmnQNJpEWkAbCnuibvwvfx2aGk1WUhFWTW7CD1AgLT1jhTV6UcxKQEn
1sh4WNPS+IZkmBWNhepYS2DdQ5vIpM4GnO6xVQcFsM5boOJMMK2kAvvkkynIW+tNOxMeMeUiTBev
62vjlEBqSdi5dUtJtc0lWe5hyNBDm7JUaURoyke4t2kXb9ulBKMOxN4rikBoWGVQZ4zx5Cw0Ih+D
06OgcYuUcJQL0Q48TLCJwUMKI49F4IY9F+bEMfcv48fUslm3MpS4BwClQ+jTA0gVcTnM9aLdozb8
NNaWI3vgJ5Yhze5spdKz0TDtmIyTxYNooG93bkURIiqn3Rf2nr8yTWRtZ5R/hyAfU4rUXHxpz4lM
ysRaJefJt1l5QhqPUn88XIawuZDB5/v8BSYLKwKsdS0rftOvVz4Ip186ddFGwnw/a6RSFl9IiiHQ
4454a7EjfTpTymTbOXGbVUlFryarif7zD+8rPEGY2z3msGfs1E95zXtWpE7x13Mfj0fYMiyyjX8I
Cw6CcL+w1/hGgAAwD56QVpQvrLcY4iKzsjq7zFkowPTKHx878ZIx0SXiu/VU+0VycLmNCAVbIncT
uXOrTuZkvdsU5sMEmKS1f05a51A2V5fePDWRrbbR3hXanofVpOukJI30qAU3EH4XFTi9PnGUVZSZ
EGq1XEF0Y16MQMQEBwCV8qhc+7GukCxKjHwwv7LM/L3fFPVwEKWqQf9v3jMN20piPKnjgRhrwfE/
ckZYbuT5q3F6cds7GzSNtLCJEwF3vKsAdbiBZ39x62tTrmFfwGuT9gt6FSNEyWLWbgwt665sJ3OB
V2vb5iJ51NLgpYTVoKh6mqXthx4BHOANoEn4dfqdXLqOX1jbYMmpNN6IHL/B5/rMpPyFol0dVL9h
mtSyrkNljuP6w/lQzHx2TiyIu37OrQ6NEGbOU2ZLazXOGJOam+oG6odKdqv0+aOR7VSo9BfBS1a3
U85kt0Bmjb3vak3gCENjEwV9q+cVDN+tH8WzhNp15+AxBBJt8MJQZL9FI4vE/6bZpvb53KnNWR4L
WjT2fU5l6rHHewc5uaQ42zhkgPwgBVsmaEMhDvlfM/4oU79AnRmAIKwcPhvGvGZlDpof8/dMYIgT
cfLxjLMuXAEGYfF9pM9aWZ5tnDwy4c+RpDQqNViMhHRi5g9DIkuEGRskWNYTGMzVHXXNg7BuGFK8
PBTXPuPVvHR7goAaFRanjZ4YcIKDdiuqK3GldvRAFCJBFRqQthsHjB0h1sG0C/8QiUFK4xYBAt+9
1lydXd38AiSp8g34fYGjLBlz7QoXeKCidVC81tFETwmvJQFIfyjrj1q/xnk3jMywgSAYPMkzzRqr
TMQwmhT1+XOQGX8vorwaZOtmn2BFO6yxt1FF8UwTEBuL+Ga/BWAjUYnpdOPYHgJQNs+HWE7Wl2Wc
jLTAdNRGY65V+Kxj/vJ8Y3uqFDyq+5AsoKl74qta2gVxQKjKTQrCIyTmQKoVQbMSBL0iZSF1+Rje
RWxXJGELTxYsZ5I/b7LcWCB0VWc8rPWjb4tkCX7thPip/sdVQCBPKqA5QssDhVxIbZMjsacrA267
IlTb7lgsNpPwHVAjmMQMLcsEzx2r5qTBAqdFy4ZUf2ZJp+llA/SozNdFqt+Dd4OHwVZrXBnQax9o
P9AYAHhw7V0XSUOzNargbL0BGFaa1yUbMmGv7dsuuf9KQgqLbzQwHoZQRbv1Wj28zu6AumR5uy9Z
gPuF4EJwqeGyR9YVulJrq/VPCfQNt3ehhE8dWFd4qIG+y4zntIfp29prCswWthFg0jfpOn/vYKXO
bgmquTwj+qhspxa0vMYlNUXgcmbuJnaqVupZFG4PulJoQO942NL2u3eoJBzc11qqlV1vuupl5jyN
ayKsLKPAxpul97Ww7MquqtRePUKUYcW0mtg6mwJg3zeGawsPQgzgA2CezKxye2CFkx72TF5I6mBT
PKmVMoawMfcCeJtLO1aV6FrTzoV8KkjUelOapm3xcKBlxHruTmPZDLxGPoG2AIJVW+ckY1sA1dip
/9C0lfu9IvnnW4fJh6ya1yUI9haXS370zDXztWjsN7eXUvg1v8EC1A2DGBcX1m3IPqR5DatfOLDK
JHBcTDtRaZMG7hTBbcCeXievD7YYDvZPFF63yTU+TgvfRCQ7IJ62LcfdYnAhjrY2o47adXQF1AW3
uBvIDpXmjjeIcRxawAth8mFZu5UbC/VG8IMBgcjNkHPHTJNIti4C2WNdvABWYJBdkS+nYvghHS3z
Hv4/rN029CPM+l/8uKQXaJPGzFmAzRPJ4nr8Ta4l3OjsYEq/9Ctz9IpQMCI/EplJtzt4DkK+VY6E
b+fJrfx6W7JlN2Nu3VBJt5fi3drnFYDJQThZ+DC3UOb8uXEDF4uq22euYvXHc9OL0d/BqsjGHd7S
oMQWaRnVjnv3RggZL+1aHZktWiKhOx6v5euhgS0gmgPN05AMnc4o57vspZwBTVi0MMoBIXdbN1lY
pP1DeqM/dSWDc0t6bT9s6ZEF/cwMsPw19ZfNBLZNF1IqaG4W8AL4RKfxReByHcxrgdjqNVk8Ug5g
K5plx8L7Xd/mIMivF4tuLxu8n2Mo0J5jGssxx0JgP2tmOBq/YH1G9xZh2cLc2bASXs5V+hbCPS/p
rN6wZUxTJUe8L0Dx1VjqE9jw9wnhVKKB0McAxM3bO7tHf4IaIxWjG2FebUe+bsd1uw7GxvpMai6d
mvCQk9HkvLetVYpxHWerUYPZa0c8Jfn1wtc9g+WMiP/bqOQHMIGzAU2GVTa1x7oF+NycnBkepCAO
ZHruzRXUlciywOba12p2NNHOYIAxOo1HDEKawmwG+szhmizfPLW13Rn+Kr3+FniNBP6B6N8qdRcy
wfcD6Ejl29espSd4tuq8DpYm0rONL+66xoexOQBOLKQRcsvDHLqXJBAp4iEwbiEcMKezY+MdRswu
uiKTod3miZ+zOPIAktrl
`pragma protect end_protected
