// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bqvmBnveO5JVHmKzYwNmW4OxTAcmIHlRpMhtx8VjZLCP0vtmbbxzWGWPeFEkACqEydAdWsC0gOiH
z+uEtyXHRDecenDolq/ZLtRK8FHMwFATaYaqh7cLmQHh32s8B4Erd4XfGzDG3QrFEUxVIqAuChE/
obLdLxkDjeEQqjy7QdLqSdoogOglTtBkB4OU8ixobC8HMDrTG4rKgk2rWzoJYZxc0kjiB1MbqucO
HTC77PA1h7I7yfdl64yDRsW+Sp6fheDS37en+rB1HlR1MxbH+eFKVu17lZk3T5ezuo/g9yQV5k+q
qKk4+LswFVxf1XHl3uSuz2i+f+5YJxDabzCYmw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
smy9rI71WeUxCD4V9I6Zw7Kv4GXzTXmjQ+4JCFH9itqdThhS6no/Gwzou9IFVu6toLBJZDkZ9cuB
DL/FhOnLjNzxMi7gv0AkkQMiNkH+WlGeGjqSosDQx9yX1xCiShUz867ATkOi4WxuafJ81sb8BzH2
Zbhwn4dtFrQe1rQw3qELuyJ119LJRg8C8dufAazLNJw44cnqk4dxGgwuo1wy1bK3Bf+9LVkId/Y0
PGPhX68rpVKya/Nb3GkQ6nGKu977tMaLScd5tFuPlcwp2iX6nfIOjIZ0EHEMvnP2xCMhsUFdfaD3
/j4nun6qwMtOHi8nlEzDSQ/VisT8eR52YnsASBx9vQaiiWcHssNvp33ErVZDqhfo0XiKuNXvu7Pv
rmc2kEmlPD1t3rH0xlm41WjSoNY0kxryVLyfWKmFGPi6t35coi5yCqiCMqPT72Hv+yDm9Blg5lDW
+c6ZM9z/AxJ5AWAPCJdLln8wDuzFIwZ7cI0H5NpK77Qfp7V6uXAEz5PsnuNqKcFmcMdcKxQTCU/J
mt4mGxsixRyXAHr29bb2nBxr5BmCv0sp/v57EVchvXX4wyDw1D6v+Upt5kOcCBDnxtFmz5kAGsTb
kIzX58raFOoj1ARrDzl1uArwy0TIMFaTYiJU4qpVemJ/5xLhtmFf6U3kRUY9pz6yK7JSJXxQPRWw
SH4HnUREYaYclpFR0fV03rs6wZOGgiihTATbkKiL98LyIhOvgwSEJbnD8BsoX8R27msJewlDkUzQ
5xxjAeYcK+Vw9iu8oESARHa90Il36NEG2Y9xuVYgOBJlvv4LtHaZk0b9h2gsGGaBK4wlQRjtnE9E
wV18bLaPuUbVG3eNX89cNduC36TlTGeoCCZf66IfliBlyByTavT3J5S/hbLPP1XEuGG6UkKchpWs
80Ui7qdjvczJWriErePAzAlnZcGC/M9u+yflGCQl40JijT7viPf7URMbYN4lf5LMx1Rpe5fXYhQt
HzR4o/EU54WxdlqV8CaqLi8gJU6uQxepuAlX+PfsrJa/fh0rGRC+9xpYQj9lJyPDlsgdGdrR3AHQ
MHwj4ZZPcR7jSI+3SW4x9uw+ceQP1vehUGlj5Ir3NomVn8XHJkvJw1qc2h/wNtdYfvZ4lLE60Ai6
Pl8tJc3VwxixkX4QXjUX15fYpo5yfr08iKoRrNvnPwN4Q7hxrPYTAn02LIJgYnf2nL44G0RW1Rgi
vm5kfnnG6bs81+VOAmVHeuBqiiEmmmImoW3FeONGI7MHpijHLXsUrPpViYrIvp6NPIuw6Q7EwOH7
cgfbi7F9kQYh/ifgy41F6ieQLROT36b+pUK2JZah7SPux+I8HYbtPI50g+niBOfF91ypwACvttxJ
+wqa5MgtOcOqzvgPxMxN6CAPrpHt7PN7svMIp9lxONXfqaRQSoTYKM3foAA8LgQhrqLzmovS4TB0
ZV9mycKOb4peyVDzv+Yg9tRRM1TspiSeApq6ImdqxZCvlk2eI8dfI6n0ZEZyyRcP79DwvlFA3o04
WlbkdsvFeCBCKE20dKdY1o122ibQSuSPxacV2I+VrO6GlzwMxsJxpIKH81mtKb6W9Y++2qbgRoVv
TYD7FWycZo+XW8/Jvo3Vq9nduKvgZkWk9BFJopl2BIRW2z6zTyM1zyaDpmuPCF3AKMwLGgrHo4cS
D7h7fXe1ZGlxHQwWR85LZevfE850j4QC/w0EnudncbJ7jYq66xe8bQ7mf5xMPd2iLfQINQD1twKH
bReKgm0CVKDArJmpF14gUHDJw/+WydlfU3ooO3qKe2TsPKUVl/yHseHRzvBcfeElAqa0gECrG9bL
J/fwDsiycJKFzUfJjlSmrXB1F0CmhZf3gB/2fYrlWoQ75J+bEWZu+tshyCU/ELu6I2h1fMkL0V44
67semGtkykNU5YEIDFpzDsnMEfss//3I/0GOySvBzh5Ngk18VFN8ula17U+EgpR8pWv8s8kv3Hc9
owJKU5RU5AA5pRldCRfQtnl5Qclwtun8yJGAHYELotcamm8DJ/3l1uxklYlkn5jOwKEtXH7ecgm1
4SbARfOZJfzoMrING6PwGUzhGVVdeaupkP9fLExXNv6PUwZEXTIIaQ/D3cSKmDLqRXsKj+ym+IeM
TN747xcJqVBkOwv/EDGF2o/OM7X6+l8MHDTH9etyIvjMpzW6BKUJ31jNZf89zvhDJ59kBftfcXgi
k9WQQc1WAOm5Qjsh6psz4TgbSrTdWLerIOuU0sUbJ9zADKgkUVsyehMz7QSc2xldzOuPmyfTr9mw
HrHXuekm0apBMU2LFOI3jC3AZv+Run27lktih3rdJBUNMMxUwypGl+l9emnblsZmf1pNNCUNs/u1
L7doCjs9rZTcP15h+I193H+rMHUQHO/cpeg5qj6WAS4qbBGJQGrYARljJWf6yHMczBf8mk7p24LC
7673ZBW4U+2g6fwVCQFzwNw44UavNiqIcoFNe7VP9DWfIQDP9ulBBY7KFmfW8pQI16Dc3w/pBf+0
wtoIHVarh4rA9Tw8q4FhShQu+tNOJbErGWF+f58bGYK6GWdrfGwZ4Wr83IySd6x7SYrflaZsQpbQ
V4jjiSJ50qdUovAU+0YGfxZReqKTGVPVMbOHumdB2ohZB9BolcAHcU1YLqcuSM3FGKJJ8ItMtrY9
QL0rLo7b0WSwNs1cb2cL2LyuqGt9sSq3RaX+9Th0El7crpYjJEqEdahKnLYrn679bedoqoo3ZxSj
wF4UBLRhNy75bndQGUgdKLvQMmKxp7ugdwnmKdpGt3P2akQbt6uQY+pXe+/A4v5NQaPrY5z/uzej
wUK5rat+B/Mq2bRVcoaB2yiRzS1kczsh4qSBXgCEMg6rCOBB6VkDKb606dP4cTnEuV5Iij6DH6WW
PD2d+00q7V6kGYq3/mMdgdrU9jGlmDdDwEvoX9g3YVcEdwdM+VLTt22eDMgz9GWxaPIjkRYET2T/
eN8wZs3y7qH/YxN7P0tJyJpU7j3lx/mzTdJ8vQ8fdTkALlhk0Ct+Mn0zPO37L2b519qNjUR38raY
hioxKcJYNxSE5w5nm8NPnX87exoTo8Wq4g4ysuNX+WBTwqnuqGtZcN/fOjBhjU349ai+6CBPMDiS
hw3rwWmEwzHeBySY7mAY32aLh5V7EUbmnT32bgCVpnBq6wsBvWmBnJuo+QmbnUOqaROpJoh8it1w
hk850Db3sDizIT9GcEC4LCAQPOC9spfV2rIs2kQpsd5QsiK+LrO7w13qVw+wpGB3Qp4K4coCoLAO
eJ0L3b0I28KbfTbPu+HJlMxXM1BGTdCXrzgkE4+wTcPoKFuYDg9G9JaDqeP81LVGCGdLDB+drg7a
ApaX4XL0knaZzF/KIXSZcQXHLf7fTTIuDdMKr7O6hjR/2VPSI9Cw8Se7v7bWijc9VYetJ6pyj4ke
vaQl6HE0x+J/ovy8ndmNZY0ZeVi5RVA1OtW6QOwKswOVNZ+xuu8BdA+2MsVJEgDzf9zSUfkkb51G
JtHgkiNGQdXNdPmC6G5BBJuXDh1O0ZgZylc226wkdBtnCFf9h8Rsr/alqNSX+9C//opFCrz8Eq2v
UC6qfOqfPcxQp6+ZeR9dwxqp3ydhqIHyKvwrSclraanTA+Zzk2kFt5/WBZvqGIlOdJLB5Lo9A61q
Uk3ffQHhY2JC4EFtYXCVAyb7UBVDZS8131sP/rZbFR0oAAsPon4NlmQxXOnrclcdY3MQsq2Fjmzy
ppYFLTIsObpiVlky9KkV3j6AvT4+PwKOK+N7PzsAugzPjQzSuVfzDpFQfcs9XfEKgRnKykKr5wsz
BFw97bSMH+1I1j3ULD2t1H9/XkuKUIpDeZelj009SjCUBFqlLhNadpZs02JU10/krQohCCbLed81
FsCWEyd8JQOtK0KoJzH+qLuHFth3RNwX1D140rZm6cBKw73KFek2pJN1f1HnZzRLew7ky00u7jv0
Ry4Vf0X+h1bkkQg9cf/QHJbFFGtfjb30j9EIuQnewq/RLN4fUdlJCuPyIEmpafZjYgRSRaCPauXW
8xlfV8BcEFlBlIYn1bAZpOmQ6dwlD5kHxQqr9ZsVetLh358Gp8at8hRO1UjfwhcCSwvNFHApL43H
s32dk+ygERUMGRuNicH7Uyt15TmebkptSTwGnHmAqCpBwPZvRqVJD8MOU4ZbLvrAyZ2tu84yM0zA
H9kFRQNsF5YOujvlK7BCebj9ZdGpZh4Gk4NDBBwY/J06piChkPZs9z0U/PqO+o8W2iGRH2HAOrQe
p5dBSzyV3u2YsCRN96ulEufTg7coZFAvyiYkCTWmIQQDN2fP7cuYMQG8BTk/DwRcpU07CQlOey4m
bhlBAUhoP0E5XkF9dmkoJSw4hCxF3w5vtFrykNa+FfOiLMkUp8NPq+ZUC04f21Eo4NtlUnALwA0k
BurtsIK/AVlSfBFM4tFzLl9rmgUqGyisj15dTPNlIX70+ralaD+mCmv8TOrfZPg5ZzqH4e7yRiRT
pTCNLebF5kzcSDwWKmzbD1fKLuU7OLaJAG4eK/zg3bJkcqQ7v2wSO/7Anp5VaxxSAmodaq8xckh9
NbDWG08YCSBhVKI3qWqiMJUYSMjhoCYateSTbiVt50o9WDwtpnh4bE0jwNIEyOCdjcyFUD8IYzht
R4/+rZCnma4bIrfMXJSpTw8Muf5o33tQeeuYA/sNoWJm5kAnky+7Ex77mAKbE6p7/JE3ayLBr3pZ
Izdag8Mk9Vv7nPChXBvnZLjxiPREGe6hTY4BihE15V6gt2qsxTr368qH9LJRQXHmnSX3hHYe3Ig+
t14n7/faaZKFGQSmq20cFaFnv85WNVk5We+nF3jPRmjFBRI2L4Xp6fUuczNJ0TmuHlRG0P5mx4A9
p0A8Ml94JRX+a51dQUhYeWJIhEG1xPoKlRrbNJGmX/ZSG03dIv/PXQD7MJwVTp6wWuV6Ztk0DTb7
gMUsRkPSTcmdSamqZpBWca+QVbjMwTigfWseQlP/bXFOAGBmWTOMlJcQBbQ62V+GwH8WbSi5qSlX
CFvo1L7MFUZ5vS8mXnwG5j8zX/ahEMd9SGSsSH+NdQp24BUspEvIxPPm4rvobCALS+Ug0jUX1ZoT
jYBVE0dzt/uyb6LGjfpjCXdvr2GiqzrrymHWyXz8gPnJHmj6Dvcm7xkjkIiyJ1VRZTHuOEs=
`pragma protect end_protected
