// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
sfRqNL8tTmNhohnKESRfEQW0f3vWbTqQyRR2XAeNBYqQMXrGwi+CBsp/6flptnos5g9aIs6mt/hR
BnDKrtQUkL1+4/QtlhiwsWeDeevyXakf10lOCpkKodGvvNKo7kr+4WdAl7y2JeNMjF5EkmJGsCUz
aT3+O2ceL6cnosPsU5/ZmmYn9W5Ay1Gjs1jksrwsnbik6kcdQoG32t4A6QeKXaVCprmRccU4iMko
UoHLxtUwZinvjVsjR1tO2bfxmTk6vO1NfgDjWfVjWghNs8ywRRbKMAimfEvt5hTtqAuicMLF/Tup
U9KAGoyU1WfreOqJ1Yceah2UkRYFnoFD7NBLeQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
P+daf2aeLndsOzqnt80n49SILQlG/8He4aVoOldAPJhgGiab6K4dDX8VKvVnQZM6bCM8ysj1eNOY
Zso36YLBa4seCloAlBGk6jHXzEfiYN6MxQRsxq7h9evCwUzhgJZEru6Tuy3O7RdA1/Qyt0VGu5hj
nPKzaKB2R5CmgjXDozBM0oMaVfgGLZ2kpUePge5bsqjbedmH4jDV0DCAUkOTzd2YBDs7Xt7lkVGW
2ERVTgyBaj2SVe+Uiw7hMrkn7lyAuKT9iuXqJgDGfN2aMqDE6uNxSkj1qp7IqiYoBjzbvT0UNdyR
S/7FwTnQTMMJBx+FIibfpZHv0IwN1lOKXg6a8j9SivPDRHe7bFG0hoKBRGh7/UuBwgvwkRBRw1dD
Fx2fPbb6+q4f8KT6KvGbuOgKq1RMcEHXUqBwkI5fw6eFaZMkW38KQWKjS0FJ5TVnGHlU7fOm8rLH
dpFfhtoj1qVtWNPy2Kp6dOybrdwux/OsGMcKATjZ9fwFYWfg3LHqAySrqhaEqCpE7NoPBDI/MIED
r+pJHOZFhaw8c9OPszdsPxETiCL3VBQBRNJxXGwVtW4sxxIp+w9lSpJJF8sIN1wUbNQeSFQBC6lQ
QUUu2NLlQtUGpQnrv/1MFSbbKXCWs7ljFtb4RPSLewyKKUMRBRIk+2519NgDQ8MCqLgouw9kgmY/
W/a6eZAeUGm9TEJoeGj+WKzc5YUfgrgpBPtahsFC5Re4GdwkBZ7B640eJfutkdzHQGjsYItj1dgM
YRicKe+py2bZPN0j3W9ojYsr7HHuWH0mL9FcwCr7jXovc5sqWBkAyTSTNwQeivWU0+T1IpxkxHYM
F92bXQbB/6nuP3wEPwo57jJBHBGqsXyuSFuuTB14iMg+FneGQkVEY5+5ZD+4NFG6brkPPImhk7Pa
Hbu9/Wnnexm5KGDdkW6v7mGGeC/ySNa6A5pA/SYOBJmMKcYvQA5wtAXra8KNk7cV8kFsSJiVrZuj
UOP5E6EJDAxghFjjiKbaPoMzj27wDsemE9gQb+X2/XR8V5dWCg0WIdwGFuKCpH/byXMpWIHt9r5L
pP2wQcGihvHr65T9qx2N/IuSmF2pvMphYarJ0ck0T9vG0UCiHzRalrTqO0gIUobNwy3LzvZetgBp
WH0Ahrf18Vja+EAI6f93+H6VKoyF06UOmwF/0LdeGwlsLahJEJsOmtcDO/O4AHyIzgTVBkqbt5IC
hCst+gjBLBiziYi/60vtJa/ZHnnnzZYSbH+fQml4wuwaZ5aa4TbYfRi4JhMKwbp/dC82gLj/OPFy
dJjOejlX5MuabA6oKeLcIhFBycjdIjq8jROWygsyoba7h+r77EDtOArjmdQ1OUWjf4K6ezzpNFcr
8Kba4xzQj3Z2iBp43+nP75PAmaXTS8g49rxI8oZjlEbnieHULJ3zm5eq+JwuXkAzWdJ09som+4s3
TzpMa3u0wJqWDicNrWU97WSSvT0MI0KHOCd1b6EONMB6a+RjhHkyfdLsngNu/jtGuZq8nTHEoE0C
izncsaYmJIrCHVIhKz4yFsSHy3nQ/2VmAdUKnjsB/hyFaPZToLsSzI3fUIeHLMqPZ8co9UqmhSg+
EW1bX9pxfqFWKETaFTXtrLbaI9B9tZMRoXOwBNcJEthE6bocAjMVMwCMEjY6799JVVf3owX74zzP
sqLi2gXIgveewFSm2ULhxSqHsVwC+V9Iw0LYr4xvUkZQFwxJcsQp1zax/hnN7/WXkGUOjoRqC0qe
ofuGNgDhoFQqS7+s0HS5cXmobU35B1OMwVuItyaSTJAjzl/UQnDL/hjzYvfkD4PYwn0PrPmqS9nP
JQ9rA+ochFuFmjss/tAb/6TneJmdtOeFxtlzspx7TeMyE112Rp8St7nWLB1BY9ORogpv7fjJhRMu
Z9x8amBPuk6RNmPkh8O4Jdg7OcrOtWrSpX5bTg9klBgPRtp4BvTt0vxrL0YAxpP5pRcYHuWgII2G
CtG/NlnmaMVEMKIYwBhhEf20cW9OlxrAkF05YgMBbaGWkd5+K6bceEdv21xREZYy5T0pr/rebCdi
/ph33zXs1hy7DOOpYoDF7dkcePoJPM7h8tD868FedGTgOtTvHBpXU6Fx67Ewl12hZfD6EheUTNhA
xkbwaeXar9/oPajnyfOJ9U8tysN1+dtrspNjsjaMmJRrHu3AIBsUt9gK1jR61yQk4HMfQ4KmRVoT
3rUPuYr27Oxhf8q84yzYc86yjjdblOFcnvcKksAji8H5YRIZDzPVIVuyP1CUqdN+WDkgcgI9/CPN
w8PM1E6rvDfkejIu51+CMnSM6vNcbVYTt/q4YTFb2eVE153bIfjNSgOzSmPNG/itizYWZRj0OCsa
L7EypPW9rBj2YOpDSY2A7aH7Wmo9n5p9K5cpJlNgQoN7+Pe0/3Hz17JFsHXBRGVwbVBMzpK8qzba
3DBZyUOAgX/kqmT05g3hqDJhlY6rdWoKE5OCQMTRmLvJdz/hThaYhllF6K1rFxSoe5tUOjmaHyU4
IZvX+JsB2Fbgc/qaaYk0C304FNXNbRARa/RXaEmktunQ1nCh1dWuy8nLjBfUDOSOYSxzw5V9FiL8
CvgGYrLPuQDi0BHkKhLpcDhfyleL+B0HWDork3z+bBGlKFNSy4huIHG3J5Do5f1Lr5vbhxOlDoJT
hLOPR0pwlwtucRALUaZSoLjPR8D0K7NwxLI+MriSO63jFhVcIM6i9rRuEi0uhzEj2OmMIivwTte9
0DBQSguWraV/xFxSZTtBbQnpuNt9RTdLzU7mLpwmSlqMKeZIQBmlI/d4Wptp2lSKQRvAo+lq5r7h
JochbVR9v5pPH4nC4XE/CZeEWhHW/gvvSIfYJ9t1wbKtbWFA/2CBNHhH9eJ7avFd7n61/WoSOp1T
9K0K/EINeSgsZDKAeQNx2O9Qbz6Wx875WbuoWws4uL9spxNrVZFWL4D5jUc1iwg7WXiRplcHyFpd
PLNdTNWbHJJEtjQMGQ6KtW0YYgaVAsv3kg/i1ZY5Hgi5kWmW0ecSeiycwWwhQumUe/lnU5RY1PgJ
nBsvbYQtv5F8bk3t7iGlG2LL7fJOVpqUe/PS+hryy4cLKU4v8veFNVhZsKAaRWOGwunMM1o7xxY9
392RR5ceMTVLs7EQhHqtTP61n3MsdMdh/wLN8KIbKVjvn6i5Sfp/E/JA8+YVObrG/AlAyPXLxtR/
wm5xHpCZNBbA82QZ2+nOn1CSzTy/ahnkosmeJerof8FTH3o75/rKYsoUWcD+VPvzLrpPU/qfP4N5
9nEnG0OCWcbzZpfU8IyNL61/P/sfNiQc/andWrrdganQTmu83Ot+KVS2gqcexUt5Vj0dW38t8MIc
CZK9+pjXHrkQ7/KaCY+DYM9njZ9NhLwgd/zNImxGT5JZHkl4O9y2T3jnkyRy0VmreB9gUh4+IqoK
kk3nEsM0ToK8gKdj0JYwmeuiYxXrx3mZkiVIgYq3Sjl5gFcW9OeGRiMv8XtzKlQM9l3QXckjD+lY
Il68Advh/upM5WfxYK43evEWOSY9ir1wR+Q+KDjDz0RXAD/CdahyYKQrV80DyUYcM2/zeBi3FA6o
/gt4LhQci/4WhEsS5ZInemhhxD82CplNDO6YfpYsQOo8ocwMOKYCGm11RhRts8p38fl5slP6kO5f
7u68U3guqIHzjBOsyUxoDXE7eI+39GkaWNYDBmU6ba/C1Yhq+2VURKD1a7I2zslNM3X/8FqgbXhm
lp4JMNsCvmDNCFKZZ1M0ncaNpeFtX6HppXnLeO8H9b+LL/m/dw3N0Om4XDqKwDwZQ4GnNrBam3Hw
2NRuNbQit2qQnC7VamypXjBkTXvHn/qFoIpbrlg4tT7kfO2sVNEg39eqTTu9Ql2QU+JIh386aUYq
2D3bIZdyoqT2LkIstFJ3rlOZecSzpmE/KeHyCvJVyMm6Ti3B9TvK3keYlbyN2VArNqPi/Je/Ehnx
tgfa5iAvtyBqELCOYIDavE8NOU3mIhDofK9PGR04WrcpC9JZL9D+lCRn0cKblqGUZeZ7UvhlwnBZ
8X7o8aUHc3nrYhXyhGgQVdOM4PQPnqZhgha2fQaCD8bjmcTMZvLQWxxo9EfNx2ulcsXxGa0ISjNL
LDcEP1NUDPZd2+XpGB1FfpOMt22BBPsTqbMTlp09QhlQeCTITW9p/cMc8f6pAZ9DIXB1qXa0Rfvz
7KbIeHd5wQ2qvNUKC9V2JNjCckltT6NnncPhHIcs8a6KSnqC42CZp2p4UfnNLVk7ma5CEOq3KJI+
UTG2L3bJU2QIBS2zghiiXTJZmhGjkiEMAD6RquhxjlnYWOgBybIEINuD2uEFvV/SbF/JhULNf50B
AWP70ZXleyM59gdCM5lSGzFIHqZX/1MbClmKO/MlkKP3QRnHlzIDNcbAaYTyeWyLqbmQSAff0+KC
bm6riPU7SdbHVoRPoUpMTBusamBXN2dkXNK0mcdhLTB624aIXFbWZ/ynhM3ANbFfcFRo7OfNR7DD
cXMmr+0b01Qvr6wKiGa0odaaoUD/6CmGpvCJLWzBBiN40Idln91z8GmywT7QLXCwffojgDJCQnS0
M+XAu9AU803oYuNuYiMjt8VRBu+I1X9ImIVXRJo3pRpYae/hoVeGLqHvygOk3YJQkOPXDVOPX5kT
62YMqWuixcuS26DhHJmCAgGiMNfROgHa7rqrvd9PZh58TwgNrDWcG4C/5mMMk17KKpONaM3f1OeZ
Zw4VsaHLurBDnFBwgAMU5ReS+ZMKXAYBgC98ULvRofAlxkiWBFdEsR+9ouF1DMga4yE0IPgdZFQl
8IsF1qIrsL6GSaQGDeepeyDCntcDtaf29QdJKEMyZ2ohMdZ5j3Z6aKuyKfzUQwm4eZ/a3ywob8fF
nx+IpsmRHU5SkDPnjN2HOcE1loh7q2GdDWWJx8JTjSFb7NjbECLPgryha0Bdpc2Hz7D50Ftp1sjs
zO4K0pLeGY6PkRX726UEddviclFMKZBngA3IeD2rf9ZprauI0cC9ynTlYzyO0Ibqk05qxkihn/Hl
GVIrt1z07LKPZIugs0o06zDW6w0W0P7HRl3Od1UQaA4XTFYY5kyL2hxkd+ikHlCEeUzbkguncnHI
foX43jG1DAgdRhBy19nB7mqixb5VFnX6nIb55hdbm7BdhJ8ZutCTLofGRHDM3Vxfy1c8H9G4KOnb
9aKKT2YEtDKJy9MujBfbRGKoMScY02hR2EjcL1Smg8J8Xaw/1ygYjaieVlmFm/t5Sye2sgqVCeqd
pZBOaNbP9Dt3TgU+tKx85Dh7owsj0PnKqtwVT+eLKHnxITG+e8FMUE8iN2aSFxuqVNp+eVeRmMWl
iuVf+w6YrrTzoyBZd1nqmpu3gdQk9yX3TEJtKWcZlSVZnEV7AiPEpvXSucsfoShUxc8p7eZ011dN
qBLAwgJe8uWh/DuOUHvP8vpRDIO9TdYl1ZBTuKCpCpvxvitQcfIJj4hNtqFtJ8A4DB5FiK+Ludgj
/GXOWu8DsRDSylI8vPrVD9ibvDSZUjpAzzSflvKjizWezJzvM+9t+S2M2PvWHFqLoVF8zodJFsqp
N6Vtpk/ujMdojpS79as+ZiJqdLLdHDnVae5Jq1lS1Z268pL4a3iU4pOv0gpWquOXd7wU9AAPnSGl
4JQCOjddsbHTUoNCgcrhTGYyqi7xYvenhmZQi2cmVvziPobBsOz/FiHW0HbsRo23I5AOtHrIGszY
Pl2tu9CZfALHvuRS4EJ9llhcR68mBt9UE1orGDZYgLuqkZoYQ+LSTE500bOY9LbbhNx9R+TWDo/Z
om7aImEPJL2PvVbWEjIldCvY6LCG0K7A1DembJwyjlsrT+2gWwcE8r3y11ZGO2Suc2M7Oi11D3Qi
h8xCZyREdrJ2q66jCJ3V8T560PCmd9AMgJOvUU4uazZQdb0RxpwN/pWc/j0YlDXTwxpME8ylhy9P
XH0t9+qksR772lvqwcXzmwnZNe3wQZnMybyTy0G8QaCWmeQc15gA6huHkFJzazf5R7+R/AGkFDfm
5qLWylt8ss0aKxtoVe90WJAka4lFp8ML2alv14Sob2Equz3ZEEdL+Z9ZVh5Ct9MpQ7ehXUwAPjoQ
GC+vOJTIY9Cq4+r7MWkVTKXCLA9JsWOP7KxinV59moDMUVLCgwOFGphcSmgToVzc79IRBO55NPNE
vKeb5GAjDIHL75F3NISgiKiP7gNJ7ttHwmv/2U/EjS5sDu10nRLlDGN79XKsR3taOn+eq6D8Rb2T
69Jn6ZtV1eDLLTrZjWFeK5DKEP4OO3soWMmDep79hPEuME1xcoixudNDfUOLJfvLAQyrHsCNdv+/
vN3KJry7+UlBb+fHFnlw88+P7lV9WqsTse4aI2jppSYii5ylB4rRUsa4slo9xy2sF2OEKdIf4gMa
wKWI56Is4E+XaPA4Exk2yp93k9TcPBUu9mzE+6olNJdCP2Z54AncQqGGPNu0i2lqYxFJ33JUUoIK
0CGYvDka7s479KsQOHURS6ydQTjl3tHJcjjiSZaSoC3cXRGzNqUUUb9Jqir5xJFiH1QcZvbUi3Fe
ndADKjU0euUX6pVy6TWbnqXc70ti5aQCRciMkg4WopS76zDxOXpv99/K48V5tQTUKSQwfbCIUcGz
Rk/BdzZul/fJ17ZfSyr4FXQmuIFMhNQg8INabi+T6VCSY4ja0Ub4YCWUDVw6LUTaYEK1syrTAYad
mF8AAblcZ+ykC0YGGVBMsyjFU1o5HfEHvxGwNdqnLSy37JJXS2sku3AB4dP/d6vMLWorGY9LPhXm
XeRZHh8tY0oSr8O7061mn/siDgc5OyEVEgjlwjLR0olkUCVYYoDGCvA+6K7ZhYAff/YegVqQK3Jp
Ouocli8PPIYPtjvVVWTkd/FfWcAMVjtXHfyaxuEHUQ3uV2eE9E0x/eqFNNsevF0Teh7GJZWMzXDc
qJYo+dqDr8IuOvc7F/WX/YR7hYi4NQPelwxpUvfIG/V/RXKwr1iWC3hmMYdOq6aQqqHQN4SAvgCB
JZ0hq+BpQu5dKM9Bwpd89qt+RAEjSZ2xlc2ARoTpJwgLucy2SPTOlVnYWCkjR9TQOxzie431DTxZ
jrdzDVB5myUS/1hML83f94prt88xpxIuACSuZqUFryvSN+BcA05zhE5QK/6PniCVhcgV1O6O0qKx
lehvJkZ267X3yHWX1q4dtPC5jtv7MpoCAfpfaHmd6ITY/SrjvgfPDqT6zaJz42ZiENa+lOxgixNB
9WkQI3ElhY7VtERI5vScsE2QtdFkVEFWsv8S9F2jk/Xo8Z303cal0JbjRgENlyPoKsM7s+X9xWfs
c3Tt7go1bLUoW2jlElA2sR+S21kZdbqDVWg+VyET9A6KjyJSd+zGGPOuqTvByJrYcKj2G1fJYkW2
j6RgGtA2tthcKqE10XrG8HBJxX1/6xodCnWl2H3ing5PyGlsYKRnl8mhlOfx9n9B0glM1nQmZKcr
PElB0+JuRKXlwpiTXie/UokqcBc4EOoUtptiyy/sCw0Smqb/xOy28SmD8r8DBV/RNOgIay1Fprpc
4VqEjUkaWFEOIF3JZmADuWaegVyGdaQRruY81Hm4rOhs2HBKuNo2Y8U7i6oLOVO48CAoaYmIGxrf
TIGxOKKxkgn4QHRgssKSHfNAgbznmaucJCamVLhwjP9t6MwrZJqADDk7TBpXdBsnLc++hDhkvJAe
aSY3c+NQz3FOoASLqBEtSeGKtnKUpDkptgxyPl6TaR1+EereVdMEbNfAX2Sv6MZgpxzgKmb77Tdn
OqP6wgjvS6eAJVFqoNhg4E4s015t1NUASddKdQD3HvLOmPe8f9nF+sDeGCsQP9CRTOAQw5GbplKj
lG/4JiQw6vuSvcHhLu9bwORhD9o/gMLQKfdSBLdNf+Vb0eb2VSAy6U7UZZSYmb/NLEkjN6xTwhMC
Eb5e2G/MKI5ftj2yodV6BLxT4hj2MhKnZv9LSAizfjC9+BgOB8O174j1dKtDpwaTdWJisDb/O9i0
0RCxZYwRBy1MxK0irqHvqZWatezliNlz2Rb/F1fGDPTsW71W+akf4rbqybZ6fCodsdvRrb1p+OeQ
o4g3an5g3Qf1mztp2ejgfGJ1/bBQsLBjPfnMQqlpsB1JEPi2u80z/O/pQ6KBFLuRsJXe3baLctQd
DsmcL+h/fgW0ApL18i7bkQcC3NoqNkzQclSP2Fog+Ka5gSqhOTv16EsTIeBUZm4gUsAsNcefXTe3
ZQO/Pl7dPjzhl91ShQXQTrEe64IvJCvFog/GgHos/RyJTWSpag9ikx1sBF9CpKfBQUpk6445Q8pT
6+Jdl1qQ7L0Qck39Wa3hcT9F6WKuQnbdw4TBFntjqjSGWhG2tuzTVJYxWWi3/KI7rHO2cyK2FdZb
vzzqfFL5wwTeOraGk+iiIhu8O01O9WQeqCy7+ao1a3IuxC4s+Y+vY1PKxL2D2HhHjTWKBLLCvzVO
XuVe3aQd8rZrhs1VSX1eLA+Yw3G6QHVk3VbJ9gzCTRlkrSBI1mRfRZttwamfhzxRWKP2dL+p+Vi7
X7E5fzaegseLwiaiJFjB4Y/Hym+wIawTBfnlojMHeazLEQGPy0crXWN7ET3Q/1DidC0qEhGP2T2V
VSagEsVmp3DCguzPotOM4CZ+3TMZNL8UqDdqpinyQQe7etPyXJFPEDV7yG6Vn3hW7u8Bamdhan7/
orrC5OOK01fJzGBf8gL6x+5O5r2r4kI1C49iptygXkY342z5d5bEyuYh8k5uKxu+stPVmolow8jE
ckfchCaVbJC9pEqZL5AKSxeHbooT/P+TOEe2q66kh+PMRKS4G1HUmI5iQ2A9sVg6xj6Raqe41U/E
KIfHMnE8XNeDCrMOpOC1i2Tzp8/g/yo0pEKlt6KNF8yRFD+vL4/rjxkte07ho/lLiEWo3GLe/Geh
gNNEN7jqUQ02E4qsa2lethslkCp9ZhFEnD5yIFxqVD1ZjQRd5iRS4boVwp1qB98ffxOdkTuBHdb2
W4K9by0CUZF44DGCA7JDWfJ6mbASJnoLbfOFJM4yRJEAVvnh+74JhhJ2qWU+S9V5JKKeHJSIhS5Z
bWm+04uvkN8OJ/+46P/Cjqkt82MaCIuO+MGpxF6POpgS90DEXr6iBmR2vFD3c1YURNCQBh0LYSes
5jV1tqOqhESDi8LU0ju5dvb3iMwTjXxPB+RsM+DW0EUNzzqaZJbPvKyU6KYn0nouZuTt0XW0D5Sn
N2sIueHckwQTzfFJKeTU/AyxUksANG9129QvSErrM658E6U9P7XK9WCTpfrfzfHeT9fdY81exJI/
gLUxKQ2dfymdzbHAv3R4YrhsZwhmzMzYMJrQJwW4ZZ6isWH6WxbbBjHyi0JahG3Egqye9dRtwrt7
zTudLQWbsi9vIJi4Jx0TkfAHAqHq9Jhpq+vdCYxFvTWNkj11zvgxQmNOkEecPm9eveOLBo53i++3
QqmVeH9G8zi/vPXEwtSXpJvuyzUeqGJc7m16egbaAwfho/TFSqXn9SWZmIUdxczMiQG8LoDnPlGX
SNGtZZ+stn4MQat7HF0mDsRtirOU7lQUNJFuBsqkEHuX9ECfYjMYS2vOfzUkxfMg/jr9Qrwp8XTD
sVVMqIuVcZAtKFu5ETdtvLE2hvp0GU7sXF/8sHlKgM6xGQ/fj8hHl5BCL/sdrvZGlVONi0a+UXIk
lD+ug1x/HaQbtpQlQXlEQbpOxB8aZni4G3XFpWFvFyU9vOfrO9t0c/RtojRcCVE/bjUdGcVzOXF2
zxpsAcaR+nOuxQ9m9ijaCC49/XY0BBrvgLNNm059N6bANur9HYjMRad36Djx+NeChHa51UEwLwPs
nUw8VuJuxe4paye4XLq58GRQe5/T+PVVOpszF2sM38/Rl04HDUeRRDuvmywOLFoVl7h+QS2t21k7
WYYhOmY5Y5gcrXF4UPgZrkQT9fxLmycJqFgWPzXdtnm2NgZezhbECaLNLnmJLz4hN2kXzJbQlONz
0OM/jtdMWBpuahSYOa/pVdF/p188et/BvO8IotyFe+uMCbYbinUyjjtK/5pEBPNv+9nnVVxXEBq0
MPcDBXnaaA4YfEkIfeaSQRRs2WTBewxTtuq4Zj0JtfPx/axNSSfEXesQ00vctgwuf4biZPF+2gZt
kHiRXasaoE9HuHz2S77F6GzZYsLYVzO14f3TIF3T/6aexJRN5I9hfjtOUuvyDgewp8UWskuD8Myf
E703umCQXxdSKUbO9UmSxe1ezWFMh2542VyuWLaXL2HT6HW74VFw+8aM5LU3jSterhBNp4f60AXG
kC8JSQoyNGF/foDk1twhQ9C85Us8J716gHkxIoDiV2pN5oalIGKOilYPccrZFKNcaPYHWJlAtOhX
ZgBsumbJJcRRwdSNJy42th5fLsNiNiOKrczNh22wDdB9+IuTdeGNijRsM8jmtTB9qfYodgarctXq
GIVWUj5ggW1hOuYgyYecVTZAzbk16ZluEAkmOI96PMqTZhFLda0xjh63WllTq7ehAGJ1qp5bzwRV
frhUjrSR3rwt6JpUqR0ccnGSjHfhMzBbvrAQDmx62hIRxSdIF1Lji6HhHkCqkt7h74PeHu+nUBYQ
CwPO6LMmk74RhyMuFrzBvZzcLcRkreK83aKV8bWDZSQGYwcIL+Ec5QqgIZhHjxA0rBkXtq1JJ/gO
8xOknX4E/OMuWbeJl5OmXr6mPe79wUe+jGgkiX+Dx7SfN0EUljs290owJ669HlrCBH57KfTv0yEW
qTixEEfNQ9K2F6Ih2/l0V3XqFK+3bCvDrkG0ojujfFf+jg7sJhhpt6iix6BWg4VYFGDxpd0+iw/g
k2PSVzuTYDc58Z152no7VT/KE40VsjzPKyMS91jbTvXeSzQ3oM3a2b3gk/qPKfeAfvg4A0EcUW7n
tWH+Fo1KT6iOt0hjZ3pSNOu1kh3j3c4fxKug2napU/zImSSmQAfuja9i9s3wmiTh6GLBoUQrRJUZ
dfHhroG+fwcGuHedUD+fMVwVE8YoMzNOAtnCd7l6WhQ9Bm4jXytBzbqqMgNSXp7NkfrLWbrJMNM7
pEyfQwkVM3eaGK1mW89fTkwWwNISPNyWC4aoZWJK7xdSH7HihlJ0fh3KJpUBbkM8KfO2qbGUEyDX
cG/uA+b4Znnj/xVrPF1m+9YtS9WKrI4Zk7z78Er37I2Y4rgHdzpqukcLNK7TlkSUNTN+0hm5It7e
qjDU8LswqxkoHbl0I3EXCgONrWbSCnGWoq0uNHwpr0jaPgtFBjmogdyWfeutfPrLq5GqOY2PZWrH
aSDarJVt9a3ihWZUiyKDwdPRtj9GI2MlFiML02W6AasaU9utwFntj69IgKXybqF/Oh01D8EKruNS
Eu3CawwFyFuceYedCeQ/46XJ9AFcnAgRCFydJQESX/3omJM5dda5pBD12pl91ZG5x8v5Beq7IHmy
8ofmfdxGpY0+YQzIItKUAMxzuyO+HuwmsqbdJ2Noq20TXl0XMCWEfhogFg1bW17Sa3/iLxbO7JSr
Qf82nGMooBuzhIz+NYP/zgGWwFEe8T39Lw5Zi7cr+nbA/06dcMSxSmJwE8zrRdIGmNWfBdEdSUI0
/2lxKCjQYcrc5THS9XoT91MrDAK3vkCDjIUnUMfRN4M96jXW84UrPzvv4qFi7yklQDAB+D25t1JP
hXyKnxuESUEEU8yMJWeA0VUnQkDXYugc7YOXlrtEhecVC9FIM+YPeLoraxx80pCu4JnBScNgVbFI
2+kcLq4spDwRsk8nzPAXOmrKMEf4yTncPJOND54jJRrQRRC1l1o/DkfAbZDXpAUjmmUvdR2u5RO+
S/6RAOyPWxVNvAN3u/mouEvilw45h/yMiKyWsJ788TwO0GphOVw33IXPzEhdZ8hXueX3aTjhOkWH
TRC+aZJiL7RpBFGRThZJyuG0WdD/6GVPqugxzLmfRjn2kI/a7JFZTGUWenFJxAEmwt9xKd8AFdzR
fAQUFgDYRG+UvQJe+HhjfImAiurcBT7rVDKUDFYG3iDZliHDUgWvhOYqsKtvaNh4daAT7zJDj28V
owYNLwG5jdZYJBS251ZShAPU4LsGfraiwcIhe7DgUNp9TV+w5Mjb0bFRiXbNqA5ot16+vQey0PZU
HHg7fmU7zaC9iBumle/N0ZlYd4hCuH0agiYYlNnotmQJrY/TPibKR3A/GY8Er8l87dBd4yrhl+qF
F7uKbFh3QVtc1+NNgZ4MO1FUL24h8vQmwm1O2Ohvs7iZUZTJC03nS8KL1zsJxA5T6iq4KvrpiZBG
jHsomMnEim6w9mpzZOl02HKt8DuK0fXcQrlXG9un9DBDPExZM5X9iF0CEUQ70PdgQTrJfVcWCIda
Ko9enc1XLEBAQRc1wJwALwm41FGEX8da/XZaBP3qoq1FCRjXx2nRvftB8XGNkFqM33lMEBOZKo4j
HnNCoHVWP1Y/cHXU3N01opNfhkLqfKAcGCbDYHvXXE7oRzF72N1Dp0c+J+m8fC4GLuKCdfJww+er
wYV0G8i65TFy1vhXIAQZ7n2SeUSv2FU8zy3QmNPbZjyi5BpalWCIOwwdnkV5HD6PqbdLLUeT8twV
Z749uhx1XZLUs68WWltERxO8Qh6wZjVTlr0vcDVRUcBk+PMeUlyhXWmNq5o6TNJ7jOUw5SKwE3ys
cPFB9MpvRwmBoETYyzKUpKVEtqA/cJE02aOSo8XtYLIKoLWLyBQcMy8+O/a2qfwQ8DEcZj07fnNT
CUTg72GdhCiX3Q5Fh0qFUANHOxrIJg60Dn8HymfPzH7kh5xbyOHl0VzV+kw+d1elSmXsSqZBb+eN
YHDEXGCWU1YwRQyHNHQDaJeJtBYUDBxiyd4dKpKZWXZNNJfOWyAHP7gqV7PMf8KclPZ/uQ56Gf3W
9W6nw0Mah6/3N4zgMDPxuPUErWzJIBZx+M2NHl+qENv3BtdqwVY9gG6k8lmvf2K1x0btptFkGT5e
987DLdC7NHcQSqThIgjsNkBP3JKTJQ/KT+A/NcLvMEn4xJ8nMPp2rXOIhWmEnfdjaG4XpJDbMxjF
Bj2NH3MYwDMZma5Gbj9aTO2JSqT0yBGaMqo1ndHeO3gmz24Zp3qL/8Apg7w8MP8OjcZcCwM1PHSj
UiwkQJbTy+IF+2QbXxotQvOtSs6950ic06/n6ldavifJ+fjfNAZ9bb/4oFh/P7VlavvEgyp9wevo
DxaA41wVEIgxCpFe6DN/Dg/00gQTLzRL3P88gfXYPusqUOPt4YVpu29QvAh39zZZ0n6XC+lVAaK0
6hrqAUWu2IOZlTyT+ssta8OKZ2psQDLqAhMsQ052uwWJogy87mTTKHXUV0Htv0vmx1Qq+osh4jzd
GWkwthrX16vCVPhC/JAwTidGg6dhi3H+4makSVzyZxLi38BWY+23M4PrmX83jSr+AspsxvNPeqi+
6HyzCcyzNWoc3bdZCPghU73nlPn3B1QeXkFXUCSgrpoKikUNHoXuRYUEmBXikh00m6tCYk7JVx3x
x8unhbqtSHi6PunmjxIWd4vBbIDE6jef+Csfvye0DeSlrAB6nvA2UmWajN7pK8uh+sFCu9mHal2J
cHfVz3cTXavmRjp3y090Pd4guqZ9JeD9+1PmFMPTXaM6Pk4YCR9lYKUAqf3qrIVoCBs8XHBp3jNm
DYpVtIS5FcD98tFX+4dmewOI1a8Fv5y8cTlKqth+vn7cKXXERC3gEezd1DKxMIQl0rgzowQOh+qD
M410sZViK549D0dVHuHnrm4IqNOUTxD1YY5yplcKumSOo98AIfhpBcVqAlziHbzQKIrpAR/OQ9b1
2h1jAAq4qIxcpuUlrcnxpefjhjvNYC78BmaPn1hl5JvbYdL1WmnVqms3slxR3Ka7O6Jf+kTso4HQ
GpSXsVRvGBaKVVhztZN+BL+it8evnYEdFXK9BcTmzhWzuXtq95yjp+dqo9h4ODUGIZcRGIJ/8eSP
tCiuqI2RtNPUvL1sjV6THomc51LX7K9YmDz7x8tJnCGEiW4zM7ggcHW4nykbs2HYhYwvqIx6QeVH
PIoW85VSLFO2lZMsXcLKBEVNGbS7+XJBi0z5Bwmqe/sWfxwG6SrE852Ch6aHV9tKz+CWwfu93VU0
0G+/e3xmECcUDdldKGS6DTTzM1bOFfS+YUGaKYXNo7s7wlliBbX6gO9rZZgvZICSGxJOHBZloSpi
OA6a4Bw9pD+9yyV7RiJxGybM0gTKqJmtxr0roc6fCscFnMC2pVKR4EJW1AlOyEwOr5sIl6JleoLh
yDI1/Ey37uep+Kb7XnOxjtM+KaJoOK7GK8lJV1yME8SE5uv3FBuzVWpXgU8FSz9fKszzUcohF5gy
3S+qrdgjOdqBMiEOEaOqsqanbqMq46AqkEuev5Jl/86bNIruf+9V6oj+Y7NoBuP/fderaqfM9YiD
qQU9cHxHYdd++ADqZd4FQLWiWLZFca4gT3EtYgINQf4hU/HWcFIcQ+H7S5Lu48DRBxlUUKoTCHRW
HaI8CdrZVRjcos5WQqjX6JVebD4aFVRFr0cAqw7HBqm/3pX8SYRt0RhhR2J0Zqe0dX62rtSXoixT
crKyQsKCVugzzzTYnnZHuhmEmqdFPxxwiXsNrOP6OUYKG30u/N0K9VHy7VpoQWc2Y0aJYQXJdDKa
iILohEJ4qIu2nDuRldyu7Vb+HGJycCjeazuwKq87JWvDq1W5MUG3eB2VZAilT7Ex4C146vH6sjun
78u3GBckZbB3UC4Yar0ZrPhtyjmU/1RlharAnG3DBEbCWROh0r+2wxLNkDSV4bhs0PffUDjHjMDP
nrFCsnFKGK7I9KyVqRcVg9yd2E6CZTbQ5huIpK9b5PZW4SOIv6prGKA2PCO7VEfLWNljnzAluW80
gOiQTs6osoJJUcDXVlPo0q6NeH6K/lBWhMzEmhjKBJwu49EURCOU25vDnEwlNylhVkiOw7gN41HX
5onSpa2r9xzLPEvbiqaCkGSJgjQiG5ivbnLWmbfjlSuaZVhE7+ZrMt9kBiy3htNVJ9aDSmeqZxXk
EAP9+JDbldEv39x/lCXHOxIewqSwD9zBidbWiHXJUPD3KTfge/9PRGBW8w75SnQNzNabVE/wd+f+
jdVsSyzTrffcAPNK0WPftDPdrQ/fiReLJIQki8lDfB0eJMcFD9wPTfa6I49v9jHH6CnOm8LXv+i+
4W/W06APHQHe+XLyMQRmv7dxPkDfccBaqCap/+4yqOTH3E+MEISojhZ7U4K3aEvnBBf9DLE9DKsR
Dl0/C+mUq0d0Xv1yGPRdom1H+cAnjXjqWfmv1+66POFC1WV0xX+3E7qAGCLWZTm1CDBaXbpstJD8
Pb+TLTSj/F+9j4s2f5w8BZbX727No9qdNm+UR4rF+EPk4irbAcrfuWoQ6syEjgdfWDYbFNvRIyDd
JpdQkxnZcs0Tr+in4mz0KV94+3RD4GNkzkuTi/LA9jD0BJwm8FPGoaeknXOsdrApAUCcx370ex6F
qVPTmjJKD7ErPsTPyJ5V3D2xIeT6L9tjTSw8zSbqehWAOnXXd7+ZlyK0g/D9Ectezf/IS12R0C7D
A48AL0RKYU34Z0ik4GXL84eudU/vQljH/0vj/cXMePajpQILneQKCWYEihquCwgdjEprJw24Eefj
+s6UmTvtpFFWUH1CReSHwdfrcHQ5psodFQAMi76ySez+VkTSEQOFXRgj+myDQ9UvHMCyCUO0oDAE
79dX1YlMs+LglaXG0Ve7dm/Y2U7dCOMWu1vXuH9FhRw3fHLevHbxTHAvq5bmrK43DUVEPvLlwjcs
zWNSZ8vqCRvq1bYyV23pwnmTuJK0LsOvbErnAoz58PbLq+0MNRkzq6n/86ZDri7mmDzCOKDZrq93
qBlZnCU8oOqaJ+Hsg3dhjCS4YvP+wiUqDZFqkx/OeCF8u5bxK4gc4Jvs4Qwb9xVR2MhjvfVqDfih
4O8nmOdyf0RUTh/WfBu/EZT5p4a/OfZC1iHQvkRl63meOxAbqemIgDGNnj65YOIhCmS1A+m2Avbf
GdceO9WO3Jt42O2CRmGPrt7VD3BE2h1YJFoETKKYNztrNOkXdzKXpP+852JoADBQC3C0r7EuKh0x
mNkJy15Ai0yUzude9JPPXkKVKiRvlKG1aR1UHNwwz+XKys+NyPGpHG8CwBK4sBlzB5du3ZOMroz8
QziaLrFEBTDJO0PtDhj+vTwmUULE3FF6tzETyJs/08rV2YgZuvublgBliJWpDQpVfNbFBv4PSBY3
ZJ7W+5Q8KxyjTT703PBnL+TjPzyWme0PIyK817/FnygznSxU4xFYUjPHm2ab5FtX3r4Bk6tzZwaL
u4lDR41fAykbfH04RMyW6cVse3686NxC14kDUEhUdyiMjvU1cWBwrj2DYIJEcW2SHvcoVrAPRawJ
CkO80WAri0N5U4akC3DtKc5RcOev8N+W24MIvh0Su58Wr2IkNkyOjo0dcPssp5PiaSwMhYxrShJv
R8pk0dkmToO2VCnJ4TMH6ooGd8JVOj9T2PqTrXxWxa4KqmH/UfUs8DjDtUJ3q9LG9TkzKfPGHtmn
fflUl90aYRfzs+T9MS52osCl97HPXBKwx4E6NjYqOlRbEDay8T5nciSvXsB5rbn7m7huL5ekmCmJ
vMmjX39AuW+1NYZZZ5yH5lXyvO2ng6StqTBAPuStC2X/YjzUUNCfxqwOWcoRQOJGvLwc4WPLij17
ms2m2OK0A8g/P2ohyPqlAZ76b5CXziIOdbmqAJaThQiMINMpRAGIgMLrsuk+lVBZfNjnISrFLaHy
ZYyyid3KpTG1IsFXhTZs/0BWLWeq/cOXGfFflXZbOcnAtAKhe+wqJyU+YWhy9COh6dcJVBQTpdjB
kU4/UbUU0ACrC+LPN/TKJSS5GnGhdw3N3IJpiOJZ1j4M6M63m7bgCfj/7QtDhIhjmsqJxqPL9PkB
rCEowy/fbQpZvHED45b2ONBkd9fadog7us2pTm31qXFX8+H5wflY8hUUZxVWpUt0Zv1q80UFrWzr
FkjAnc5kkrWqLdsEvsJJvfJTwoQ5COnI4I0e/WESRezbJjRLqsTCI+FYK2bBpREM9floles5oqKi
TPZMRoSkAmKGA9vBnBTXmFTzpAROUnmQ0e1hnaiwiENDtzsJ85/Hr+P4pw+DhiQoHqy1nNZBAQAJ
1ZuewBqKTTKq8/2OdGGdmquYCfWAjEiwdzTVwaH4yjhwv5ubipbLRF5yvEKisuliRYddti4TZvAj
98GZpqlAoiW0Q1COYfI4jGzFcu0cVV7CfCwvLOBprMtg7lZI75GOxDZMOJ5jPro3Ax8M6xoDI1FB
sxortPhLe8iOBMKIObjTgCYmhlpK8pHHHahEWIr7MMM0zdA4yCh8yJkcNGH7CLUUGGDYMGX3jiaM
Vhwn4qFPengh/2kj/u55k6Xf5tmiPzSkJmgLYpTG2qtTJFaMv/kSEWG5cZ3G1JjdxdOMq5m0s3HB
MzVKWLBEF/4/GYPWi8tW7N1c8pTwSfCs5Z2V+ACa6P6+FPYgor8JsP37UwsS38iHLCa5C0oqrTqM
DKgtgVcDWSpBOgJZguOcXQyPADThQZOltjhqxI2lQP0V1kiM0z2V3m8EuR7fBUb8Ur4quuRo9Fam
nspvMtOKFoNp9jUWyKxIjXgsNhVVNlYTucWhOZslhAkSO7LgquOpNqweUg1zIm/jUabkTqiX33ME
XytK7CeAroQVNZkM3RyXjKsuxthz7JyZA84DXqsYaYZfy/4TfYlNavYighQCWwzBTnRXXYYTZHBz
fN3VnxuvidFDb08c6GTdl37ZIhkQKTm2glP2yS8W2G4pxYzE2r7WSPj6mNNx1LBJoYwtrHoSJIv4
XZs41dwiDE/5oWN6VeRBo2vdDuNV81OWXTkfFL09DuZ8XQQQcRpBtL9MvzrCwiVqrt4RvWIsfscX
wCWNKvZZSrDwSrGs2d6bBBr7T6R8im/bC6aiLjXBC+/e4GH+zJjtfIioowtWm4ETVkUsaBEUc2PY
WUY0KdDC+ajMcrp3W2vaF8F4VBwE8CijufTVSAHZKaguBcjZ7D6daqdX/lIXaC6aV+k5t1EcatNs
dGhHZj7F8cIb9rR1sSMs6zuj6CFHlGAVqZy3SEvw6E+aL/M++wrQ2uf/t1Pnmma/x7liNn/zceYD
2ljqRUgdKgdOY2F2sRklVyki8RaY77eX0ATFx2JXJxzo7IQqWJ06elsNsp/g/47dPZSRzvrO6Sav
TDUZgf06OKvTQqfLP5PF4KAdWCpArCmucrM29XpqTJAmauAOskT8U9hqo72ykvjvvJApXUaH+ebk
hk+LaAnocZ1tKGCkho9QYBD/p6UJ8s2QdeYPrfZRwE5w+3GejlF4hb5YC7KjWZo0kUanp9S2m+Tv
eECrJHm5k7DhKcC6gq2alxdmA1IORQjhFZSxx4jvozE+iTgt+l4j6qt1J7IFBpmO9rFzvZp3hBnK
0BL62P+0B06Np1vYWoQZ5SULtj4rV83kXAIklTkw4QoSsJOmo06iZt0uYqHPo/iwpzVHEdzxgCEY
EDUK3AoqWaceotf/2pz/NraPVs0Xmymp6R5xrxlC+LDsMYqeucL91mvvyw1BpaYA5XwIm9KXRM4v
l0o7jIL5OTCER+jHqgHWJSDiO0EVmmLbFphaepp3rZR16HpOSfzBpsMUx22kswf0j3gjKskCEGsB
3n1DMMnnZUf14lz6LMexYcMKIRJusTw3lJBF5uby4p1Bd6TFrWbjnodP87CTLHB5+20gzrUExteU
Nw71vkamZkrf/4C8O4hELB1jsQDKlLkO2GAb6JTjkG3Bhi59qwckeatwU32z0LD86RBKQhbE/jI2
BwUm8kmyT5SWsmvjhREd1zu9tJ38I8AuNMIlvhpzuhwaoz9IHIaHt+rodLTWykaez35WhTUXnu5D
jGJeBrknN/H5tYJDmwEygunv3IewCMohjoBT7YrzsJD7kCFKCtYLukG1rgRHKzE8HoMdPiGPtzTD
r70WZ5Nj6Xmg68RyCclexzXJ3eQEgsWHX3AKpn0Ia3TQHxpDiVIdSQwc5mpJoSPlwN+kgAnUvZXR
yvn3Zp4MBhN5jokasgDSUmaDCBCIn8PV4uHQudIazh9Q+bZIToiGXayync2QSOgorE9gVCzlRnof
iz0Vtju83EAQnkQRtciJvnRgRJ5Ih0WnpPaskeefhmP0mkaRqHxMR5QRgluVPWdJ4LfoPEB5uFl3
aK6iFgVRS40OkvcYJeno8jblbvD6wBlvFDhLvX8a3Se+AN4NlILfPi4jRd267L1aI43YmMfOc8GA
KrinPaDw1n65yMLkzuipgH6Moba9ZjbatPt3zFSHa/18RpojuhBgqjAoCMZam1LZOaTklqH0B0VZ
/EwtfAyv95vfAD6XXyK4ksbcD3D8qBGSQR4DAz6MHT94zbz4HswFX/u4lAby9/YQ8NuhIlFWnXGd
bIAO9TgFrZEtVMUvySAG9wuFGJk7KLTQqRcLdz68bC3c9XhmKCKL6FeG2kwrW29Xy3Mg1aG9uxDo
GdB4hqI39QCU6JmresjRwBuPWdtu/GyOF20ZoN6rnbHdM9Ez0uvbCaTwou+RKRAn/V2yYwDVLmMj
8Pw5yx0MlljzgZk54g5LXiUnfPgNCsaGMn98I7CFzPdwnMRds9Kz1LTivKfnZfdNx8R7jL6iVIb/
1jvDR7ttZzXxJDhsdx0SnP6Jdh+eXPKzCejpPtF85ZxloWMKc2/wWk7sORx9FRvvaCyTSyD7lSDa
4W4kcokwQkJhwFG4T7sq+7Z8y3mm1ROFTjklD1QSST8ZDeVtZahQ33vMxnq3EchVXm8U7XrSHnIy
AHLtFwG8Ewbpn9IrjAtPvIMF19/ItWmHGkKyiOu2nwr0d6bdQQ+5ediArlu5QBvZ1mPebB6O3imZ
3Ux/j2T3VMYmA8aXzBJrcisapxzq7Ir8WQ6VQ1nFVejQF+g3gIMJ1kHTXLsAYEiwCMjkuDhG1CRa
m8oe82bfso+oNJRKuD0c2d9noL/sNWuPaMQyYALyArIj0/IhSU8yfQIOHDxZf6pu6pE658PFCz5u
ShTzh2DVgC5e4v7u37tZ3E7ZkihxhB9Oad2s3e2PZQNn2lCWM5zb+qav5TV9Fs9a3hEyla/LZd2V
eeQlsk3C8MBUDqk5CvRUs9auCXCpgS+wnnISDmBJIPkm9TJrWc8vviZhPheaiM+ZU8WGXhSwevZZ
b6iXqXnIXEdk4bRh9t0P0xuqHZyWR+SIzeDA6BFo/sw5X0SSwHg9E6ny4P2eCC/5SMkx9FIdryIc
pBNGO7vKC6v0i+fECFw6r8Lg2HYpZ6iRaQiix5uXazjEVdZtXUBGWk6xss2mq0xwhiIdXvGycjAu
xMmRLsED9697dOe9Gc0S6gZk8zMPGoysJst5qfNVoE/SubW5me6VmoaWIp4XjAW5xawQqAJ4a2fm
4L4dpZkM38bqku96RyeS/Ik0za4zPG8rrVJ0jygX9H+YLoilvjtQW40t4uCa751/6rLzcdyI3c67
TxnYXdHKz8A1yCkGs3Il1fkpjDeQczJqgCygQCCQ7DD5ErJgVMI4U/RyGLvP3iI/sAoIZ15Cpyh0
YTiUebRdXpEJ5vrgFPGnJTJOibVUqrZiU1iZCcpERysC8GMxHiEu23zaTUTCL14rBZXwyHpTwt8S
1FNWGwLgHj6C3r6aGJRr/iZ1QgFAnKFhsZd5Nk1/Qju2poU72RpPpxklkWCyT6gY/ELrpGf6igra
CmdCxu+jueN+X2hNarFjbDC4C6huKFs9e2tV/6wwKCNvJd7m+1cqN5+idjwrH0lSvzedqm6uLmy2
J2qj1GYMVzqb1CWuZkg0KAOdbAY9qSpheKdulu+A10VPHpshjeb7PV74lgqYkanAf5Daitr0yC77
RxGIpb4CN+1aq2jyKu64hiU8WEJgMTMJVGRz434hrwGftiQIuuqgMTNo5T5J78uDtPDHcWJ6TLYy
zSbipyhcdLtkfaDxT0QJEN4Q7leTSyQl65MKhIFX6nf7FgKFJGtW+RE7q6uzjrQd3f4MQLpfkgjI
XjykZl3LPbt0A80oZ+XhEqD0li22WYxQPymEE103QEQBEkW6ISDRGXC9gNgI6Uv5SwGPidyVIdz/
VTr3Bc2bZlQQAevmfDNXv3vVorm951syIZ6KghKY8T9sBGacA8LwJuS/A2o7Ij+vxRwzOekj8QUC
5+QebBSUCcN71SlG08AygUVDkRl6AnAcmnmpEz7JH9A/hJP/2D+N8udnUI6gpbbvUqblaE8JPrHP
7JE3wF1vNAjrVMFbm2nmZqE9Lv6BMEUaTUe3B1hgB+7KM5ag8o/SvE8C5wuPsESOcFWj3BNtaDTY
ZHGS3d4TN58OylxA6/8nbJyJqljlpYusoMTbuEUa0sI8wC6WvnrHpfwZuXRDdEw3mTtfoqafXJ0v
QsndUDh9VyvChryVRy+/KRs09/BKO83K3DCOZ3vxmzDIooWksj1jhh9Op34d3DHD1fFzcBvY4h4r
l9c3da+12eEssRpoFwui2V+FsvSAfKBsp02E903lB8mXtvvbS/J7KYPRHPWvL4S7M92kVvenVw3M
dnOrw4nkPdc5U5YorBK40diS+PFeIEuIlXBhRYPSgbOPo5M7bfb4Ujm2QG77xeB1sVv/IhVq5KiA
HIWcbTzDSAa1mlfBGVc6UXSp7euTsO/aQqsg4AR9IeG43ZlLOHfqfmYoEWVrmyFhv5bVRsB32Idx
NLRr2mS68E6Et83zVCgIPaA7ervBxQwLFOSXc2xRHorkHwSV8abmxLOrlqcv5QRCc+A23VH/b7eJ
bCZIgWdwiyAvDwoHah2EC+ubellf/cbFyMFi7w6WW4TPCWgEnINJIEQy248s+APdPKrN4urt6WcG
sf4PfgiJ6a11VwqGdej+6ey87PRgUyKdw/inyMFFFtAQDKgfY9UYsF9U2KjGde55/dwuARb2uKpf
GVVuJnBffQWoWThSS5RCpv4FkDstFPgYNdTFWen2T/kPcbeqtcYA0MosmG9zyQfbZpbZ+rlv9dys
40UyURfkSsXe3Skrh9Osr9NzVVP98iYmmR0GfqLFZfw+5FgRaRDC2hU0WfRL6tmKQmEY6KmxwIRj
AoD8wJhC+YVwERNCHVkmKr4id14O6Rs9QahgMJJ5sw6NCzA1R3ftcu2TICjJrCI7Mux+C+yT7Z/7
TLWMEuqLI6j3umPX5det3S+RyCsdZAvNSu2RXkaN966QoQ4kYFihbdIidhGdDINWpGir3TTDzNgZ
WyBdCvtbu3zSjI9EB5tYSLjiux/EZcjnVDq8ATWUolLRNJz5Lpe9XBW3Gi8wKKFu7LXlXFhJUxXf
QZgvNLQYT5U4Blw25gEAFtJCBa2cs8PDg3SFDc7+R3MeL6M6BIAz+xC+v3PVHZ5kHs3EktfQMRy9
hbi/znauArKwSajZW4MGh+AauTpvmV2X4uXuL0pLrZ6/4SWSigCYShlk3rTUhr6MSmTYpeQOuY8s
ahV3wG7eUbareB7T5aWPEAr00Dy81pZkIEOCr4NtG3sB3n7bSMwnf8jqbOgGH+sSDkME5SpDRHMU
/ElDqM8MK0IPu/MNMohuEgoPMzuJo3Ibt/vKQcCmNN60k3nRRvyblM2MakCw0rF3VRcQ2oa1Mx+H
k2DqaMCS+Bj0Q7YLi0dIk2WTaGTo2k5NJYV9u7R54s7dJPEfkFI52cuIA9ZGyQhi6bI56Yxeo2rR
P+md/WAWUu6wWOFvGOVk9xqqfz+91VC/fiZQGszIcMonhpPeX6zxrlhLWebWSmo0d/wqQavNLJRw
NU4KcNNPUrEtj6ONII5SWEjmcExtV0IC4D2mf+vxmY2QdXXnmrPNNDGvNSc38gAaVEuKTYgxq1rn
tlqQMwRnhNfX5d7ZInmUK8GTlkbu28akxhmdVhtkCWiTInZSCIGZ+XkzQmGnATKjrdEU1QrejX1u
wSeQgvGdlLfS7NrlF/Cz2riN2ViklLQiB24z3WzCVkgFT6xpAcOJq+u0PSYbq5VZMAnV0hXaxGpn
uZQUnHA0nmj/g5+8a845Z4r1H2fMERiGuPJIpDo/2qb69hpJhuobOtkoOnDmnTo7A2NF+Rc0+cbg
ny0ffMOZmI2eHQF36nLOZU7vDjsmwL2U2v9Q5vj3JGvyjiqz6rNiJg4+QEP8ijiaJ9O6aLJh7Kkg
Ul/mkGlzfgYMcGIyLnZ6oMcGoJpQJU8hv4eygBK4s6knKA+KZkn0yavhrk3n3KABiuSQzzaBHaWz
ppesvVynM+SLAUeh4uITvI9CuA/FlBJE4/BQDymjUl0Y/cOfriW3vC1woQTB6uZhaxfWU9ssBbk/
3PCOdM3nMe8rQJwWpZaRjlGPL37B2jLPHmVc9MBOJkZC9uATbuj74829NI61Qt43f0hyEpkL3zXz
3w19WRUgR7ELlvGM8O4z8JFKfpS3KdRSE4z1MMJbRH2a7XgcDZmIejpc6UXH0DI35t17tUoG2+7i
woz+xgPiu/zQLSmNQ8egYKAoZ8ew85vK7wRw5OqHSowkWuYM64qvEzQ6ZzoQg8gUN0F09m0+hPGi
D4EvCdj2l80pvCe1haWIg99hS6ev+PlpwsNSpzfptUpq7q3kV2Au2MAIqVMfm8JpFI7GY+uv8/0y
Ar/FzsojhrCtay02LzLLMUp4PTn2SucwRdIpwyNrPhvtHIGmndfA0GRS9UXqHrZLnqDwlANngJNY
bbAB11eNYm9mdVaJB25jIca6c6a2+Xotazji2QuCb+B2eCuznyEAHFqiY+hFUHqLMfsIuJbf3A8Q
eSJkNcCH3YJCsCf9YYnpv3KxPiP0tn3qyu3jk5lVtbob2W4k0q/jHs34mGXmEkRl9TFyRv2FebZd
aLqn/A3PuxQCPAj7qG8u//CSmyoqQZRF5dhjl8Kx5nYmfgIc65k9/8pWngdVMVQh4+7ZCGF+4inq
i24qqtRyMoULmyThLRXzWEdrZbJfhP7WHoBX1thVmkT0B5z5fQG75Z3uPdzDRr2jPYKs6bWDPem6
kM1YVQunzS3xEh/EU3OsZ2JzNt0Kyn0NOjJl0p1rvurExZUwMXmco6472OdNJboL6hVb8Ylq7dEm
EaYItsUDnvTAMTLsTFhwHyi7pgSwnM0uhEfv4ZeO8PfGAvtGGs69xtghh+uNsdpSMAQL+rpZtEvT
KFU3BKStQ71OS/snC6gauFxJSnPITeZu1pynSmMNIqY4mndYWdfz/yDdTFJLPenBDn7c1MWYVf3Q
BJ9J72GVK/0koUggpaXupXfRB4ia5uAS2FC9q6995hfv3ccI+n4LP9nO6zE/4O5N85nccZzYFQI5
Nu+g2O3v5p4DzCBA8Jq+Ar6laXqmbW6p6jhxSr+vzw8FvdQWK8elmIPTRD3X80LgytU/RH9UN1vG
6fsnGpdM9ysJgXnAzf+RmbtBvUKo6yaZfSoiLyfVvRg030dq1SxrWa0J9p41rDa/h/46JqnUQKvw
ebbmWojCsU/BDvFCTST84SaUiQWd9dEtnZ1xuN8qIox9iYvVmFbfeVULJbbJl1He65qKC5KeVAoA
tvIX+2bmhukQ9+IJErIbbO7zkjtxWax60TFb0vRUeeDkiNAYkmTWPh7RQ4Nj36y8a6+VJ0jr1N4e
V3LZzigMvau18DixCBEChnQdBb3S541E52OtHuq9xBSwZ+s0CmL+ZXsKxKkC+kpbJe+KrcTmNqkR
rRR5sgwgp3QLgsY0ElfIDRmrisgVHKpOk+ISYs0SXeXbFD9N0Qr72gBJV1HauXdY+2AhwhLxZH64
VEamn87GwiQP729rkkyhWn/LCec0DTGNI7nA+epT85LcCJKwlMF30y26DnByHTjzlJuKrPeId6Cy
VQQ0UkCkSv/f6mgMIlKjW+Ii/yyJ8nUGTSsetCNvPcFb/FRFKcPVhGuLBpxQr2OfMfCfM170h13s
5LoF4L58RzfoiSrSZGYXXc2fptyBDAxw0RdJbGyG7hhWdr8+KdJ6nCBSdIt540PSajHbC+iFfScC
2/2kew6/A7THs6ZFOYm913+e8MsdfVckd3HbMw5bgja6oKvEXdIarOUJmED/37G9VIxqaN2P79+P
ZMkR3Kemf7Wv0xA8Wfi4clzT38+eBL3dbepwoMXNZSPIQfUtKBEFEhZQ9BGC6mfve+x+bCtX9Hqp
bg4+6g9z4c+hXEkDZMDU7jhDSFc/xQQxkNc8Bo/TaahqDdjLqvo52m2wj650CA8YhZ/EidoWZo8p
O9jDcB6B7MNkcqdnuzvTtTKqMrUuQQVOshB96W5821kYY1zYTO0hrLxdQHnCPZAjynBce3DWshiU
necEXNRqd5WAEf8IfFYxGE2+Yxe2PesT7qhC/Tr+vuATTGb20RyfqSlnZUE5H+hLkKu/YDLaJhwV
7+JTWHUQmKY8QibL10RbLpvH/xkBdNoADA+/l7kJTb9ZuNE0flYF8gN7Tk1JF7OEVgF8hOWv9ML2
DBMh6pq4iBAxxYd+sNB6h/wIjizz9ko/Qxtl8uh7B2nJm5sbsLi7AK6yU06w7HsloWWx9HEO8Lyh
/U0QlbnoTrDCee9udjB3iKiYEKWKYFtIzQcmW3e+iYZaG6ZyZPo5XlNGnacFr1DPVdctKEjoN6fX
dqEySurYnuArtaTPXb5Etnqm2dkakoGNSMq1cj/rInx/oyASPGnqTYLQU7rTfdet3oQ4OvWqlOYA
hIrPQsoPNzM3hHGCUB5a70Zw88QTUJ9KRTUuAp/8WTmZ9RCrV3/lhoylzHzsN3FfcFOSmBQIQVcV
F3d1RxETaHWcQP4NGXkAY+2E5QXC1waBqXDFrL+c4qB0VwsooU+Sj6iQ01WgtVqDOLgva9XBjH3b
LkMoEK4gJOo3+F9RJsAy8zzjwHuQjjdq1KPUXbFPhDEC/pqYA15A4w9zZpxzPUXaAC+CMB6JEs4q
Yrf4ci6MH6OdFxWZSJdN6bG9v+itDI/kVZeshDGVyWwHpYJRBEF43MzqXWw/zoUPTi4B/yv9gobZ
3+D45x7filRsEmfZm1nvqoJKh47BKSHLQqac7aLznP3HICprNwAZKpxcv+CveB/dQ+6ZdnEUTNZg
VUoVNMYc66duYnOIio8A0ia/RqLJg1lGQ/EMHN36roA0TOw1lOVa5SiGeyIN+P9GTv39TcIEJkKe
VgUNwGFS4Mg98E6DeuDJeNw4WVi7O9J/cPWZGITEQXSz/yQ/KfpDTicRODWiDW2A9exLP6XpuBsj
6Bl88Hl0ZHPHxqzkmnKqP1wHzvr8rJ8EPUjjKXcK8i4EHfGCyvA0DRlpFMDO7OJOn+PlgFax79pw
jpgP1W12w6b5tjA+DKaBz6ypTy6H1P2rJdWE7zCpUIBgVcwb2ARCFukgLhb24AQ+NE3rQBvNYHGy
BV1jHLU+HwfH1QjBGdjQHqEwpjDxFkqdL1Las6T4AD24eeDZPkKcjgzY6WazOjpMbOmWIXsToi4c
9XzkZF4sxN4DXncgidgU6l++IM78OaE7Xrk5ADL1s8pQHMi9h+eEcpcV1PIL5+ebekQ5W9qNQn8E
yjqxuSIEZGnqUf/kXYMr9kcAA/dUaCtcgWyFTVKqlUtgjLai5G0BLENpUsEzCU+rmhfqIO6OYhOm
bpd59JdhKQznfyh8Q9B1UTKf3dSsWMtxQMjDnxBCSWAbOn97LTN2goV2ENc7zW3sdFmgjAtTjnGW
0JgtMingLjGgg5MvU9f4LHjO7Y6l9QLoCVKAswEDKNf05nph1C/rUWMtGZVh8Az/cdECeVQPQ73P
B4nFS5swJ2/28s5t6r0w9US+PpHWkJ4qia6fksvETTIwnoToJ/rgIbTeVyDwGcXTqkSAnYLxMGIl
432UIerY+ArHUva1cnca4AXjQ+O4xueTPTONyEiXLieBhryFd/9G7F2C+SwusEYkZ9HAW6KAZukt
hsnUsO2PbKQ7k8F7DTNJChAcnvEi5+Ib1YAZoTBnMuYgDpto1DnWhmzYXQ4Dew1ROt2QVtLn/hYk
frx0JYZnRYbmCqNQ7DnsO9akPAUAXOd1G45YpmI+47WnNPnnvibk0D7uYu+/FrV7DgYVv3nB6OW+
xs2xmYPCXBlejOZi833PeYSWOjX9F6bl/5bzmsFKexhrdDgsSz+oOt8f+xJOKwCw5pElvEMkjfiS
hf7KlTPedXwy2vaSThRgScVCXhyVgYoA7cwvoFfr2SFq13nKkSlQI9lf9YAYUYjHkhC60qtEsnHl
RnYrsv/VUsuY6LASmTraukxM6KD3Au8o8O+5xP/zx0zJhdrxqwj5D5cWXaEc570OjvDRyAM9NjDm
Tj1Z8Z1Pqhv9I/nqGnpphGDu8nJCMmB/CbF2QFy3md+bLLooXGLuXqJuYjvHG+xHGqf/evSw1C/8
S5wsKUCu47QAQScq0zTl28eiGavf0q2RHAWvy43zbTPlwSxU7Im87Ncwwcr9nK8tkiQD3g99S+f3
l/e/m/mNmkExggTFxup4SjoaCOlksSgHg5WNeh3x1gbK1qw/RLGIZYss/98jE+Y4ElVQuUzOVcPS
7YvnS3dT7QqDTfpgU2a7Og2fRn4xrDkYUxbHDGo/BPD5FLO9STUBw/vPMdwYtgOMQ4eaW+b3Jo33
8eOFZ20ukBS0EWGOYZGJG6c/oMZQqAXoUOaMu/bKH4O6Cr7TryqbtWgvu73Bs6vWCo84fuVxDcWx
OvyT7KB9ltFP3L1flIuLhjh0Y/mHCrfrojaWuQKLfuFJS5cY8PY4vDiMcDQcV9zS440M2i4gAlwS
7v5sAfJtne4pWuUh5MODceb236XB6KUwp4thWcXL/O1bfnPKrUaIrtuc9m8mMm250ezqhqaqkITP
nadxGVYpp3gfWi0cXl2+fbjqA9jIdDlkMaNJ8UB8Nv2J9Yo+gJe3vddVcIj7J7TGm7Ew9XRtxqiS
y9Gor2+qCpSCPO8P+9OpHWJX7G4QwTzbRa8PCeTeprcVhQzVrXjDgHwmciCJ7FTyZRHJgt6P8VPX
S3wYzzDz2BnCiQUZT46Agmg1pRR5jnTMsQdrZGZuvw/f66ew/KOXFaHKFWpO44ixtyJVDlxa+iKk
5+RLItDdMO3xlApwd2XaC5nyESiIkWqX7lAhbgh37E66KipE/esmm6D26L1YxkhP1ABdRYjvTRUX
V8/2tXzC8kDfjnOpyICHlQztIwMpyxePx0l+UaO4q19B3GQ3PhSwbt4meLd83ihbhZyNUkuImrot
nql/UUrXks698RzAVOQaaTekwEdoGR7SooVD7agzudfWEZaKGEGnIjmnF1lT8AnqAEYcIFqI87oA
Wp2GVStRDro+n3Syq9T1QqAF5jRtaAxG+ffN5q1FNkNWjif5KUE7RPwTSje8Mrx/tF0vwa6aaJT4
Pz+87ucv1+iS7yRjEHlMVgOC5dC7Hed9uq+ZTfbwe9DoxzxPbUdZV9xChy3DcZnDbeibbPhOVxoO
JfGDjWp1OPHSjmAVEc++OIQgrbW3YmyFXkmIJxYDVUIepxMFrjg13fi/YcmHqgO8dyvL0MDGMhrR
MHs+/NNVrcAcY17yMu8wcAfrsf4+nkFKy5G/6EPfxQWGfDge1mCZnGzoXCAprCF/zfk4j9nlXzfq
iCbcSZFCYneTV5Gm0q475TOgSAhAWffWLlllXhtfzTXutU41ugHnko89C1BPkiwCzTJruENyuDS8
tN/QHGJzx8O12VOUR4Nf3tySO0a+1yREcEoQuWUSm1NLYDpoGCJGcN9f0Z3wX9upZDqw0M4mcX4W
Woa024zDQD+J+bAmUFuBI4ulyzXOQEJ54kAmDLsH1M4S7QLkKg+2hOm7ootI8k9qD+NhW5ZpLPwf
IWA6hI1WkMTqB7ogNQ/AnQzxmGteVDc6BtfFxHL35yEgaIrlZGgpQnbLFinsmqWxOxHga1pRDrls
FppdJ7irJNOkDj0rno4dYFBU9xUB+v+u6BTND+8bAIEE6u56RSOOj5cjuFwZPNBVmaoATfnqehXz
keBBSO3xpF8Yydztz96qtg5shW74yn93Ftd/OjLfErOUYFHh7zT6av9eXqoAsGwCsnTl2zN7XtjO
MPnvx5885hsus0fk4QAU6uhWr9b390szQZdyu5DZlh33t6nj7TGo1u/DqTWD0dUopBhAw4FLUj2B
cl3gQiNyAlngRwwppblFRRFrsurtMQGxk/j7f5D/1498Bgaq6cZdCfSglTipYdjWaCK9i01KnGM9
1h8/UpWOn7gpIiurs3wpZ1wp21s4fH+UmxSS2Vyu3jRVQHD/mNUtt3h8k3Vxp8K1tZB03I0RfPjn
ET6mjPjr/I1f9/nufFDy9uEtEiLlsFqV4BoRXzhB8jIKCrQTngHfCIPHuAilyokRDnTvtJED2i49
zZZcvFzauX5Nt6J4lvaKhK2ECeragKvkrQ6CvjWyCndSZj666bSPyb25z+F8d7E/CrhFaKTJw6DV
r8MenwR/Go7udZdoQ3TkjmX0OXJnI172udTc9dzOsttvhyh2S0e+kGVbjC7v4wfwCmGpFbgW9t+P
NyYodLN+gDhwTdVFQfir1/LjB3U48JKiVXX94ZA0kI8NdXWATFi1m/QDzsWj8eE3nNCj30SDRUrd
UtgsVnGiQrDtU36y279yBUtdJcPhs8cklaHg/RqptIDeisR0YVT16+6rwQdOBL0Y3+Tk/IC1DgwJ
2xt2pK2PV7nMVhGa+ALYoKNyXQy0IbgTfWagIXyrEsg93h8SeaeYfygMk9a8wnUWzO4nH17gPEsB
2Fbr7y4uX9m8EmHPx5zvnOg/nB222sMumGJ9uIeCRX2UwHx3fN9qOHDYF+iVzd+sPVgVFBAdzOSt
npc4G8+wH0l8RVbd8UF/YIUWaYGfLONSyHBcW6WnkR/NMOtx/FWIbbw6MVh7+YZqp0XQDr8HiBvI
m+lnjevVFmMzV2XROWthi8W0a+gzN3quR1jMw7DD2dmpWAF0G06OUlzfKeizVESVsJDKN+dm736E
rS6b5EfvP0yg1ShhyGmAklk7Fs+lCa8mlbamKpC+BqORe3rdYAtLvKgkLDNR4VhZ4Xr+yEpTHPvJ
BPH6RKpMUBK9ZNkIqPGAKLdeNGx+GkBNOevQ792VkxPLBE7zx0UNBDrYuSIBo6aLClSvtpVj7XAX
5/w/Tof+LmAFEJn80A9uuxt4GdtURnwNUtbIKUoUSsd0AABq3rGm136ID7PCgXaFndlUdHC+Xvm9
BNl2NiPjm5jBlUVPnFxyYwXiuZUK0OruTN7MRnyXb1g4+VIEIPI7XQmZ2AozmYrsGTJu/K1onq0R
/B8qLfvxPs3w6deZpm12ha7Is+dEpSdHHHxbuHI2KZf9pnPNv86qiZFYsqqlnFfJ/SlDtK4GOrEU
dr/L1ey6coe/+YgUgfqmDvIxPsSxNMjGdS2MoUYTExiOMgt0Rb1QtjimSRb6XnDfCGwDD3XhWAz7
jHS3avQkiOR8ArWLZHdYuAk7i3DKbf2o6rg2kIt2WZ6DJflG7wy3zKsas7PMimxtX0Z4PIIxRYIk
PPb8Wgwc87FjpyCYyWZxMhXw5naTBH7+19G0h9D/9gtSncnAv4o2FskwNUl3cGQ3SmolCK3prRC2
FOvLchR9J2id5y/TD48UnM5CADvpS7ToyFuieLFFoY26hYBBhROIKcKdwli8uDJlE/yDf101jC9S
3T6MSTZVbWVaTBYuHJleB59zpOFEkhMmCVoUUogKaWZRG+WP+2DJpBM9jf1gggecZD95GiRyi+qI
q8uQBcXgrCH3SlyQx62SsrZhkwXjP36mfiTxl4fT8ZBaNf3jggAA4doD5g4XDPIHaTIPgu+5FZJM
imVJFt7bOG+rgph00uYE42Gx229aLO4RKQ3ZV5YPPF/Pt7QzdxzHfyujGflQFcCodIAFBxsxcq76
049ZYKFd/Vvrp5nU9zn2hatBFpu0xRaLL90Akujip0r6bnCYqaL+VcngD2ol7VLzl5KyXwuJmcyy
OxGKvr54QYUXEVXI4HxwSOY517XckdNyjhYdmintpRJGNDScLDkAwvxIyCXqqWY4JponmTTnlYah
aK4DTsTviXDoD/uQW5hT/ZydlOwRX6F/WN4zwWstdT0hOTcMujwdQfT2uTS52je2W3bQaSCBlgae
RjCVsTQfgrmK7Go8uyEAVTq1GpdZdBt3Tl6wTkSwJzHinlvj0qWar/xQIdfvX5EHXjnYreUfZy/0
NmqWY7LGEomlz7LBUjbERcWheCyGbrBpDTeTvyPeSzOfRMKIX6MpO1LFARCLH+63NUC8WrU/VhRp
4kc+3i79A4SYL3eLaGGXip55FKa1xZUHc6GAkDpcdx9YUg7KCpPExc++RUgGMzvxafwi+nOwAZmg
uB588kBX+i2ydhuiWl72wfqndfBcNZjpSLK47S9z837LY6Dc6uoS2GMeDql0MlNrJKY5eQp4DFa+
LQHaGO+v9zImVPNXi2lfz8fgZ/Rw/cJ0GhGqj3oHAT3vqYWjOMomc/QTbQHAvsnKFwuhlt3ZHqZB
SCLFhcDNlWC/zoJF2ETowrmJxrxRculM5ObXvX7ndmyADGb5ShxBYtz8G0o9Xqj7Uh2Xgg8Xzrie
s/E0oOznXE7F64Z8u6WYlALVw6OkqmUn2sp+hYN/ySZgdMY9wxyDE9f1zc/4F20rZsJPU2oq1ocZ
2TbNny++kEU9OR0HCjrzMzIiVfs84YGJV5g0sZAAyZvs6RSoV08fP3+goqnsPVLhxBFmSHS3QZJQ
FUOQ9bxmHvMRmTGDiV8kWNuqOPQMDQkGdGUM0LIElSBLLN8809q27FRyX8IXfzV8EstQiE0nDGT2
f6gZdfqBqhbsm9w+tIH/3527yZX4IeqRXC1KCx6uoEufhazRFpGiVfgyBEuvTftO4EcrkrM85zQ7
FU3pC3FjZh/PwOeVghqFGuiGXv+hS0aAxH/Cf2howzAcO8lkJEg/zVV4CyW5sMtUJli7JL9yMY3y
Fr54SGbjKkYLEJOcq80WtZP9rJMoqFy/fpyH4/iDdCRCYl8pZakp5FgB3LyIw7m/WYrrmIIL90sw
BJP5dJYGUvsqliPiDF7uO3aatedo9Ciy+YzgdvEzSKD+cKXhjMWQMhtHJeXd0QVTyX0huYMg2gcs
Eb+vtT9BXDK+cHp68e7g3F5F2VU0kf4Pv7cPl5saX0ZDCk/XN7HUBiMbqfJeZE0MpFgqodo1hH1N
sp7PDJwSSRSak+H3f7b2TFk5abcinEP2QbEpxrLB4IU5Q1dbhhwO2QimFZWy+LinYK8h/DHSWMR7
FDjT+CdcrScWiIuYSrqV2knY+Va3y7aDlZCJkbmfxJT3C4hVKT4BrUumXlkpM2BKCq+rRg7dUWZv
R5onKcV66Bq0y7OAIPRTQjODDMEqEzyzqRX+v/PoWXgH6eUSy2ae1Vcd3AAseeV53HVMIls8M1U2
wxnRehZXRnNXdCffwAYQdducrDcDEVho3727TJTYWwdVl3K+usM6WABXow+tiacJ37nMy5HGvb2a
9uQ5oNZGHmqvtMYqbuSEXQMft751TQO+pKfm1p011+SqBJB504H6uXHqf426/jBSj+/TFNsFHxg/
uOQCj20R5b6/M82wDcOk25GyXqT92hgXb7HN43Q1gVVCrfqdiWO5pLwxnMl6xxYaUhCPjCPsZFOL
24BvNY55E6cb0Ce9HDZCSf8Vp2nj1+HgiZfHE8TyxS+d1GwaICprVqbNpTPpgJlrItPczxHXNBQH
OGhvYK+w3LzXYP4HScbqQyue1yXjfhDRVyvjMRZ/oJLYBWFKuqOLMtM2sXc8IrbGo6z0EOk/B6PZ
Kbx7Jl2Uq2zRj/Q+SUkmhFB+4yPfwmJ4EFAvt9LD3MqDNVfkh1P44fjwlYZ5ljmxeKkPfQ8xtyWg
QSqqMeqS5EMsm8IbtGoBo+K5Nbegq3hitLvWI5KTfPXh9MQDhvPvW6YE0p7npwLZuWcmTDe13tj7
OqSQuUlJl2krQfHSC2TnB1UP7ilkW8VdTP9pBQDi1ya4xdTKrVIib1W83gGseefGjnAh+IDobKCF
SOXAuJMqoZP3uw1/kKP3z4Szgork4/VKEnPzLFR6lx71U1LDiwt+UmqaqWMtZHdzMy5ozLPUjxf5
DOJWHXPVkzbCwWNHGvvxccmyMl8SCVz8eR0y3RSbi+O1KyfoXEyEmE/eiIlbtwyjC9b0EVTB1scy
ghaWshEco6r1mq1j4lHufaq6JCtONRl0vfyblf4o9bt69FB80f1PskWJ62mwm/ynuTwzziEA9GHr
ebJ1s8UrEp/Df0C5ubYAMAhmN8Cj0uX2pekf263Xmi3OLvEwnMOyquED7wkk0U/p6P4zJ2tWJc/Z
h/God7xiECJEhJmXraumpox8aKMb+8YJthL4OlfbtTvN0Ky+GlbMAE4aR9kCq+bAf1aP613B0GS3
4XMp1FmJ6p/fiZ9jfuxnp7pau4f2K9qX90CN/koznAf5QJESIEq+OSlVapdrrC3lY+KzoEEVM87C
YuMs3ot8rccwLKFX6vuXmqvCBlhSu+xurSSmvKslXnHz5DZC0ItQ2mruCeC2mclp+MSH8RqcsCmb
y9sfeIlI9JmKIiLVg1LpvvNI8qh0cCW+TefEoQhMXYqXXmC/kwLtqSQpaCH8Qyvm/df8Eke1nlml
l2jMQm1RewhtgE6XwHvHtITPCf51JvGcCB6vMJm8+2mDAznu1qtlU3aS6ypotGkLRmK4CQ0zYQZa
4fONkDdSNYflPm3+Rki4DVJ8e2Q67r3b4IwETSNQWE+aeurgelN5VKTHFGBNAV0fefMtKJzUUJIp
QX6tUXgeyrb4FJqEcoqSB4eYfFuZf/Mzg397HbxqnRTtfj2Ia40Qu95Tc6ZjuYH8c2mfgdlzQNzI
JKJ98aRz6Uz65I4WFtRE/Zrx/p9y42MGkoMuFecgUX5LKL9WNikOV5+OQW+Pw/n2RAnj1ewmg/aC
kbDCj1T9is1koO8TN6RSWiz+DXijWZmWjOArEZmbooaWCLOKUFkFML/Sb55Xu1t0M3y8aVPwhn8W
I8tApJ6Tb+f0Uuyop1Uc7knF8oGSGSGbKP4N8K3VC/zCy5321Mfa1tDhTF1QpL887UGA1FtdpbWg
XTaTQKVB6Ooyy4jKi90nCuH/xJOPl2OSVj14Rg90QxlJ+1tWwbDN4JCCMtDq8x/SCVirCVIZ7iKt
uuq1Exa9wgxeL4FikPQp0QGfnFWPGMo1tVAdEaIofyEv/4ybmD59PqYwtb35Mpi1x/L2mJbfokho
YS6AYddxv3WHTEkL06/z1kaqes4oDfDZNL4FbKCn+LcIL16app7h2Pj1kBhqbVVJYdz6cz3mDRKA
vc1Qmh657wJOYAPUXOW42OEE4RVe+WIFSM1GPoj8Hmk3e4aAPwwZ52EYIGY85Rndq7QchXnwvvPI
q3BCcl6CWpa4hxPBx3nSl8mY99uCsZFsgLvM902QOOwO6x+VBumYC1VT8aa3YEMVEl/Bc7gsQPj7
a2GFiS6PFiL68XJZ5rql3wwlzRVpZjOk/YRSuoaXhLIUN/SBzdWAA3D62EQZRVW0K9MTfktluWRZ
oveAtV5Z4a3IXCzStWW+OTkFww6UPLbVAAC8y4qKYJOgKYDUek3+u/HsxcMnQBdZS//UiVbU1kcd
F839qfbzJDnJt2mCsDfXsVN67PoiDyN/VsfwEd3S3+af2Mua05eX8JdUKBtrVmSZ/rjVAuXFB+q9
shTpeLTawMXSEp9b9x+AQU9OfFTUwUIaPA5NbdjlML/7LOd/UNUk9OI33//ndIgApAfA0XY+qBWD
2DDiwrnsxoT7QMCh9NVPB/IgVbIEm8jbU75J34t1+e6ZXmhH7pt7s2gUGFMfsA13u4i/XrY8oCLL
VS2qEEjhjUmP/4iJQXVj4JoEte2dv2vSj+n7BQkhm5XOa9gEYSHECYeLO4mcavT+PFisZwtMIZey
PZniB+KiXZxVAwHWnnuRhTIXinsOEBGLf8jbNIVMtNHi3COm33jb7UDe8+B5Ak1+8vhMoxneYGpc
lWPR0Scp7NnlmyaXDb/Q0xOtimlmRWydfImufTO51hOTXgPwQDGrRpG3SsNwzuTnR/rdQp3AEBx7
Ai+01kWxgcitihBH1kqxV6/QxuCE4m0z6Nheb8Yl3aMrYRbWL93rnMeWIFxog88ii15eU1D/89y3
O6riycjYutqCyMFw0+EI/Q2lfBZJwm9GYU6MOup8BsfOI2GHNS0k12NXWf2lNPBxG8W/CQIgkQOZ
BpkaaphXMCbmUxUe19NCb2DoZTI5iNqW+Trmvu93byWu+tDx3BSM/5140uNyANl3nFBbZcazB4/Z
Z8IC9o+lHeHvGJmsldSOehS550rCJxciqkrMajxXcsbiD9qAdBtsnEmS77w9gg8GSeR7guu57b/d
UK2FUBUBaYO6n2R2kXL0f4mJ20em7cwWiIim4uWSQ2g+ZncK6lmhxdmej+I9j8vjrkNNBuzw+ALQ
h2o5IAkRvSisYdKEh/8pti4IDMNFV13rdxA8mpWxtFDvh4G6Jg1HbmFlV6HsHDaLrcIJ4krBRiCk
pWB7ydeGZMIbUnwuTLa4m4P/jxvmPf0EHo4Xd9UYqyPhSlOg5fkqg1AsbWQn2JW86RxrB9u3PHO6
FQtoZ6J/KL2OXnB/yDI1mbMY8iMrQPzzORJFZ9RsiUTcQWJkQ+l9mLpFiVEVrvLP9yZupp7c0/at
QTT0pJRPM+IbuiPImpdnbkb9WgkWN02xbQPYQkLzrt90ueFd9P12gGbRL23yX6c+eUvhTSmtvZ2i
UQpJWWnHDfugchv14EkXm7iXkh72svGBqdnGeecRZ3jeHQX2dwr/WAPHBY0bYiRtxptvN6OE7qvD
wPMEmTyLs6/4B26m8ma9HaZJfE/MYx8JUupBg+ArdOU3YYZNjAITPKUcZJAI/eYQBifn83X8gjF9
MY9TObxoJMzafDmjdg2hurN28tIT8snylNPgst/C5TLmKPY3VHAJmnKfzHbGHg90D5H5A9Z9W93d
eGbiN08pGk2H7E405STJXoM1foT3ykMp8t+1owON7vLDQM5zvu8hAPgafFWTjfzpSnhSkJMHbFCK
Oipxejjzfg7NoPpkZ4MIWdCRaZDs85Sd/89VQ4XtT52Tw/pY8QgTftiwfFWvMvTMuf8qlhJV+vDY
aa2hBE9oW8DUMWgSTx0T0dtVWcRPV71tpzMwPL3GBY23dYg6rP1eCX3eg2FOEJ/RY+fk5NGbayh9
Jc+g9KXjKysQ1JHBVfK47u4HjNh3T4ZxxUafRoEM400pY+UBqocTaigxCXK1oPKebCrkyG/3Fhxu
BvjutwCXdgObvPmvQl2tKEO2WIi0rHhEIBrVWGLmUxn2ZCFKpYwuSZiXaaVQeH4I/Jf5CYakq4D6
GkJ6nYIDHJlaennn0zwtoi5s4ggFL6p6TN2yuXkXrVad17606P2jFbtAIKgzvva9KevmFwU0aUog
9apOXhFjRIOMEoVuEU1ZMHW9XPEx9okGBebQnvRoDE6mspaIETo58Wm7+zC4Brba/TV0HcFy5dEm
k4J7eNfzYgzLvqIhWYSl0Kyl/K1AKCNuLL3Oe+BsHo4owKi+0BJfZ6RCb1ZPSBl8cetRhSMCXQIl
EEEFv+TP0kf1snDNPSZIIJDYvlctsVfpj0gVwevj/InLdHNKDNb++uuucxqMthk8swNPsk1fyRzr
WmIyb6o3CbMcmpZ4lBhrKcz6oyFVt8jGwh2cjNErxM4eJmyTbBWxfUzzc6GspQo/kHnYDonD1IvJ
4W8uqFoWysY/pNLqwpd6cbnsuoGlaQ6qW57ajFQHzrUcUFVEE7/sH4aSBT3TF3xuCz7cPVQK6MxQ
7xFMNNmoUz15S4+IiQJLSp2274u98lK3rRoIyfF0HYmDLywCeAUCY/vbUUT2uJ7fxBqwon7HAENI
diPFFnZbq3OFBLBVM6gORkkqGwQp89ZBN0aGxNd17SC5Zuft33LQYizadQkaTgZLSF9xS878m6fY
mLLsjn09ZpfOaf9RrdLRt4xBrWhZBcRRXX4MB2uTMCPbOMlP5JtYXfeZJpC9OeVVL9uWlLG5GtG4
AeROk0QOQoURxj2OvaaS/w5HKFQqu6NyxxkPSsD8yUyAGggESt0ht0t7BfAtEw8BpX7XHLbgGUvE
GABs1BWkb85i//FlJH/NVnFxZMr/WzryCx2xDkej6cWsQ8nsiCll3zzCGr1/Kc3z7ZCddQQKN8e2
iHnifJwK8zPlBTMtHWfcoWGfjJQrPVoRdPnZkiC8JfGDwRXptI+njweZcJ9I4gFFvhF+qFIv3ezl
u0X/EBHe3wCEHFNdQMpDzfFwUJOxB7taFo0VZjpmpa9/ClwUtCDoS1ZHKLZVT0fElotpPZ4Sfwlb
/0JdWgd8fPFzxf3lHAcqPlyX/Yjntkb84/htV2arJAWaEZF++EJdU4XmoFJe6DdRAlfjlitOHqdb
kXeGB9ih4J5l2m5cczfgYqDOReEI57SGeAV4uZmL7KWFBrRmn+bsGKJLufKSh2LXLK+ow/fbjmA/
PTHaGdykbtEgdfpru+Y+Y96F6jYS7/iAGZpPUXspUZytVHFk+p9yOj91rU2bEb9QZ0KsVhyoohp/
pAsqC0nQgLbYmyGrqcK2pXMn8CoQK8O0FcaU/f/Pf9L3Dy1gn8IMnzeT3RBouPr/138N8IrrF1bz
R1YHakyU9YE33ZtQ4tcpeSNAAFGNNwqgSgZ+35ZjuukiSLmLLwPv/mMASHRCXXQ/18ic3nN935MN
UCusMBt6cLirX90S7TD7tLR1wOcyMuo3zIHfvzYvaKYa9i5EIjRJfRmA49QGtN4FW7cHXmx9ychT
nj/pAQoe2O28C+TbBiCNqc3yn51LRsa3ro3DERmnJOiDVkPkBHCJ5UF1ZcFc+ghTznplfZmOz2ov
xy5Ke5TiEDkZKj1c4MZ10B4HlCPQBm7NcVfRmNwg/j7oJiGcmoqPrzNedZUdv18ze0YmBUMehRXv
hy32ldHMWdPXbFzfynAYiyTUSmW0qL+7T3agdO837CZ4GJ09/L8yZFE+CeKZxEwl826b/BG0LlU5
4bCO388vyPvRoIKG1neXHTd8jOsQRqPBcePOaalZP7iCBHDK+oHFQRu/FMV7Lbkf/XyS0ZjatPqJ
zdAuS5g6J3WUThL3itVjMme2uXZ9YKL/oBV6pMD7BOpc7lF3GYeVTEpylzSQ0MITlpVpZkLUCLqr
U9bxG2YSV7IhBdvO38dJUu/9HOr99mOaZcXSvmZiEMGgTWRHgAWvcQKcNFjb1MA5VAP1oY9XeMOy
9scI81AqH8pt5MxPLvZFSY+A6em6Zeccp2xn2Q/fKAKlHey7A5sYGFAoGt9gls7cLq5dUbHKkL38
FR6yjjVOJW0PBu8OEucocu0z2eGKtf68bh1vOk1t2FWveZ25j+jFPXlHGVY9QxK987kuZUS/Z5VT
7RJw4j+pQ5QOicWClZS3NKNgwbnjHNWsywsVPQef+YIzQwfL3XWo67P4cbf7u7wCIr+oNs7VvGsR
PDX56zSrpb+DHyY7V8SfkerNeqZ31rn0mcc9qcq4Pa82pBVZ2X3eIvscqSAE7dEKSs8J3kmd1ZNB
8GaYIG+4GtYyve0aTTIiyg7qbaeQ3QGOr5v8VWF6cqJJjzw7ax64JHVqIBNSnK2ya5Q8r+OIp28w
ybJo+bHNHZ8MwUmyYjIh36tR4Fgcd2YpTMNVLqpqYWEhUS5ZG1M9saveKbWeWKASk2sEEs9AZ2uB
VsIu618IL8nqZzw3GrE3+U2hu+ZLwgS0Gp8DHN0R3SZqkDXLp+HL4sNqTgAUsIIQ8F2f6Hmmkgl9
veOhQW02ulyIe/4WkZO/ugIJWlA4qFwqjkcTFzD2epOI59DAZJrkiMcE3v5mfeTCftUqvKO2n380
77y+tvgcFTZ2BUEGcGbT5zjikKq5eK+hDd1uPsiQPZC8rBXe2Ng8kdGUje+WqTTYgMdCCiQNi2xB
hJmx7zSxTlBl4oIFOA8ord7pBFjIvL6HYFao7UJNuyio/gdnbSh5pR2M8mtxp4yUxY+P2xrCDGMv
FORuvVyuL8Kb2qRnCAKvVU0xhvIFRZtRGkIfeKHEvelzFpBQ9J2CZKUK3IdoiLlnW9iqn98aMB4Z
PruYhpAhdCtucJP6On3fsPYghxKPY8NLUTIpVUDbtfbE1deAR8Oe4iYs0Pauv9f1qLCLRxCqup7u
a2QbG6esfNgymmO6GAnQ4W1Q1Sfm24Yc+apfY0tzcKQIAp9HMu6QqwzWRmEMirwojCTmeWxMciCl
wpFrb4I7bX7A+AXiLGehe3Red/YUWFGFhJ9OsleU7FGn5YBvDQDnAKrlQ3bvvF4gdh2f13G7u0/d
LVmOtfL1rxX7S+2BGLBerMUv/q6AMgyhgaB5NmZu+09KqghWXAT2jg6gpbEIA/gTdIMtezOOApRf
II6cDX0P8Z6XXaMcINybdmG4kQbgIx8ez5BjGbD4Em9BgKS0Qqm/vZtuKaR9/wSxvmW4GbUv/nwu
ngTty/5uqwdPlb9KbM/2pgL386Xf9WjYLW0g8lLksMwG3CBPgQtLMYKxAwiODcbh4bkyxNTwz8WF
m1Zxt7Z03MzWWn0D3O7g8FM/NprWha3efyWNB0F2poGNcr2bgleVImsH3V3TuG/93u83wYAZpcWO
UyGc4E6xkmExSfR8X2VsAOtq410lLGcU2gzqMqLjfodgBs/yUsvxQyWgBDVQN1QHUOgK41CFddMS
sMunULD8djKsaX/QnovfjbOzDyemeru/pVNXv7EFvtM1tcbxFPiH/qEz7kOXCrivXjyGkB2zuFTr
yNKs9LGhMC2AvF1+wxsiSu1xaOPTwElkIWUL238k1IYr9+ALvZyaptIiUpiAXwJ1cckHAQcYteHg
DwUEpZocSRGWDZvsoVa8ZvWCGsmskB2+41Y8yDBOca2QwClJZYriXVUDzKRoRlaRYvidDJv6w5ld
GipSP1GtWLH7Jcr1hXuvLTXG2Iuu0vrzZW+9ZB+qqlyuDhQk7u8DxyhAZVn5XnP6uG1OJXci8mnx
/z6quMO78DQeGPLvOMCC2K804zNa9O/XeVKOtL9VPBQfoHfSLZ1Qmc2QMDQpEAXOUx7EgRsAWRIa
zDRGUXszomRE2YAjTQwp0SmK7BmPKRoX/TJnDc5/sn07R9jdjXd1rKC0FHk7OcZJgXvtyG0btqvt
VQsG/wSMU6Sc0kiN4YwpjnMSAjqGDaEtt/7VOBgdJ+QQTMZ7YoSgdJPKvm8hpnlqzHlmCf4ra/YB
qL3uJj1VSoK3fqv5SlwVpjT8azyoNMHOrpCb+rCtXHdnbU8607XVDCJF6JuQp/whPEiQS5tXyIBR
IHWwKIKtfJZ15eDE+w1TKaKK9qGFmuW+ZDOofJwSUefLqKbr4bsGI9UkOB5DwmgdUemjrHMGB8rb
yl1DP0UGLlHTB31Xs1580H9teoEsXbBJqZBiFlD5nypYKQGSXI0nPKkJHG1UQGyjwKV0xue4/g7h
XCYR8O9KAV1LNbg43ayxOMxSVLwhRzt6pgoyfQk/+Bk3bYJHe3VgSugg7BT/MVIqBYexel2hi6GD
wdXNoREqbzlWdV+JBHe3zxrRKXrYOcDcT1EjxN8CR40EDtiqIp7aqkyUXO93KXz9lAKx5lFMc3pY
TtxW3cieXxRPT/tBbGKK0+dmJdaYcDPmI1FEWDow3dE4gpyMfi5oj6vjEpk3/DqWlOgCyXiF/uSo
qmU1fvQLorb5376LNcIsIBHb+PFEg7ntePudwGqxquNupp/23aYnivGSCiYvgQekZZCc55R4Kk+g
rDYazGnUUISJX3KYbNGUsNDkJQKgvHhKv3Kt66HKQgRtc+/RDCIqO1aPOcFCtP/0HeVLIYXHZrIU
eQ8ehwi+WbjrzK/lhOdJsJ6ETMs9ylJ/T9f28pTUXgjzRo2fHf/xXh8eCjCJRmoS6tXeugZ3lrmT
CtqVJ5603Oa5YM0OPBfTt1cAPI+k/4sfX7Gi1c+VsvSo4pIaeDlwAXqYVuDXbpp89r1PP5k8Y+II
Be5+TuH0wgvrXOKW/B/RBKT7xOqpZlgx3TSmU+hYVxajwgbrPNyKjJdnXzb5zzYPGsWnayKRiFQY
cGOUT9G6UzW/Djpmo8RC47tTfv4Z6rUp5OrEzdCaHeNZD+ji9jU65SKQInlvewAHQ33weiBnjtRR
q3dVK7geIL4vZlG98LOPXcRAdNcJfmPxWmUojkkuCKA4fLuROPqkTtSXsonwFMd1fQ8KRXVkvUoX
yS8ydwgUPMuZVWCwH1hiihy5sUznAsql+PgeE23SQIjsO+Py4BtmPS6jBlvMIMqPoLjFAxz504dx
NLMTGllgpA3eiZ9d5CEJUnByHX2drTwZcK7+o9FELoPABPqwMyKj0/7fVsVo0KS4WGHY5xL4Jc/p
CAeISh8QaOjmqSSH8VDt+Fj/3IRMS5231+SCnUvdOGyl3qGGPWUIUUlVjDpCeWT9JSK+VCkbxJyg
WzyHA5CPyDVWciSJVtVHFMj1FFtq1HpTPl77jGUo8kK3MvqGkvgshayzrN8Qljr9ZESOTvknTuwT
1SQUaxnvHxLQjNcXuWYwcrkj5F87QIPG1VX783qZx5A5DeI4gkXhNmPrGP0+Hzp5FN+g99rTNtOG
bm+pketRGMwCezf19WsJ15EC4gts9hfttkJQu2vGtDZJ1SJfTRFBk2o6798EYfDUPCVl3XCeWoHy
OZNvAumTLDBSOfIgxaLOk6WEFcZc98rJuqTy14UD3Yc1esUye88FitTjigC6BX0KUhaAJeJaFnCH
iG+JPYHwleIcjLqM85WTMmV0ctGTJYA71VDY7Tfq8YIHm9oOwcgabMi+nbPUbNYWYRIAcG2G8sJ6
mDyi+12A9PPp8ew0RBdXlyasaUrkTZYVrTDtOKpzJH1zJVXskFDirCzFrU9q++5jZzPUBGgSnDZX
iXmLjKVQUOXClE+C1XH96UDriEYIJdzUSeULpmVyU6dpa3/2RGA8yFfVzwYay561dckYCXNWoSlP
mLdWIsuoxuoKFow5ONwgfwQTE4l6D0sydYqb44XZFS2rKaaoBpu5UozxNjh4CAslQ9I8ad6+BAWS
kKwLKal3z1Rz0yJ6clx9mbIwEkFoqVtw6DKVQo3IQvUyhMfQPI/ft0uXNtbbSy87x7POeid3hx/x
u+fBnrhxnGifCXz9EbkA4tj8Xf1Bd8QsL4gKLVIvDwk2HoLoOhpH0zU279GvMJ0w/8/jgf6Aaezw
IMhRyqoY6uqHP0m29NKDsZ28a1sp6RbeTsBkBS/u8ZrJCiD/5Qb8lABlY4vy1GPnTTocoy0NWIzh
LphnEBUgR0wNlg5vIvvcCka7F4upQK6dE2YQQw5Fgstsz8+jCTBMFgCVk6LvmqkNk3pGReUy1zRu
YjSKWbGSU4lMtGTXVM2qGLzMf/5qDEyduClbpKiLoRcpEoOzF3dPfX5cZUs2rMGdm7J+lB/yb1jf
FZJmzdCr5OcARAOCNn5fiurwhg0e/0IBxzSgSvsWnvaXO5vExYUPfi/3ekYrVt5tXfYTyQJ47gFw
xqHoc29VLImtfcBg/DYoqk7u17nru1T29w1K09SRMIbCNHgMFDzVfdbABUeAHUDYFzqGj+Sety2J
R6FtGMUeT5H9xJDnl7jNvfxKzk+DIxJmEw90HwUnrxSRCtNLxIWbkOvNuttTRQTTEMJPToyxELqC
OxYxUmokjeQ9XDvdKQOxTbmHCfo8NYx71aAE0KT8fdvB3/LLTy2EaHCi6xmOREFv78vV57xAExaq
CTTUGpRae/TTwEDOo9R+cyJCsh+kZcUmvXAkyc3kRMYqXCDVt86ncXFqc+ZAPA162a2N6qRl5PMu
F7SlBuzleW1W6jG5JQZRguKm1Q8jlUdEgYA6Oqcd1eRQPSdBi0FvUkAndIjO+hkVWEtUXJPXHIqF
3zPiv6IQkjXCojeO33ulDC/L0gQEmbTC3qrjPtnfzlGuQDfGQzy5/FPsW4EzwanH6drxcCTE4mt9
dLIyJarWqTuHdVucwn5k06x6QwQHiVmatsbqQUyfo92fA3olDVTO9yXFsOeZvokqL/QHnIgcmqzY
k7LGqoTuPhTW6oM+K668PjOC5dNmK5agvqC7YAa8AXBSGKU6nmIr+eg6UfA5Pvxp4lFGADjsOOHW
8VDI/L9GesmJozIkCbWL3y54S4IJfdDOEmMFnQG4XSqD7ylJfkFSF+z7rX+Wc0+PLbs/W37VxHk5
9yYYrRMTEaXqJbExTA7EkRBL1w/lZQMkZiwLSDrQjacbMTrL7j9I+qYLgIPEty0+zOOQDUM/wKFX
6dSEbuxhUk8HBq4aeLZD/WECA/bj6Jpyhk3U6JVDrrsAVjNqQgKYmbm+dBBxlJ4YlhoiaDcsltWQ
EXk5Y1oPdE3/QonXzONwyw9zwhiTJAaO/A6/vP2ChEliOh9dP2jbtytYb10yHmXGPmfCs+DzjkOX
lM4OAWy6LwMjA6W7BEn9+xHpEdR+KQHxtZx6E0vBoKklS02VTbWYJe0AjuivwHjan4dfLU7jxmmS
L+z8m/jl0zZ07NaE9yfSSS+8bsGqentZmYYqsl5cFOG7InW6W3cL2taqkI+SjfmCqLT+Ll4kLWDx
Dt0n5Z7u7VoBcIciKAA28lDafmTQAeYqioxVeNZAFQYfcSVjgv8cIO6FJBau0vxVmQbszQABjDEg
U0TJnBF8Nm4kLYj0/QUSkBO32hlbuNnrUfFqPVIvlcwH/sg+JM+DPGKMt6/mWqyge4N2xsk2dOMd
EJOe+x5F27OZjXVOskjFpUW8dAnPFJqNbCJHFzf0weEMC57AW5bO4p1gmJccFjdKoiJ0WvIJY8uV
3xYU5hqmYu7YbkDxvDT+ed1XkHzq9DXgv84h24piUGQBL5o9MkATL+8uvlrLVNiOglgLO6vjXLQP
5hUqX9cKKbZLnjt3SL3AeUFBq2H7uNkFbGwTsuq4ZtkBxRlIrpYsDRXTfibSme0+wxD+PIwKmac6
P4cBaJa4v5qsYInz1xBffUe40N5wGXTes2dv5+2pgP8eWMop42/x+42oPkFMpxRnNwAnGyFp5LPY
qgHx1u2gPPMgx+LGHN4kpAERyKsWp/IjSgb2zO261VxvpHCSmkfDlCMgbmNYzeyBLeYO0WDel/FP
9werJC4qSiYfBplmdLPXwJZIxKgk18lOwg8eyAO6gC8BhbzIGbwQZNYSVUK7Kb82s75SmygkwrPQ
hPm9+M8wgpEWR334ACzf0gl5qIOqXlGOf5Tb0pzRH7ni5VVSP+QAuqlWMDdFpJECRA5wWah7QFIe
RpHxvVttqFcNA3IfILiCjHdE/pm9MgL2Wl6f/psXzXCAUtNJihQoJ0mzRCBBFsGMBwXbLxIh3zcT
sc7rxUzS/CLE/EpdbnLlB/oCLAg/T5AMT27Hp45nrtEYX9hfIxRC13aOnNFL+yb5dm9v2UqgFcIz
0S4C8rZlNo9fEligb/KO/Ne1bOOfa0jsBVYLHs/00mlqO9SPZj/LopfH+LETedZISPlwS+eSMW/E
DbECm+42dQiJrmMIM25qs3g0rfBcWeGpmTAto+35ZLjXZEcu0hMP/zSONzxJjpftMHZny9MDunCO
0FQr6L5ppZ976FIePe7LpQOsODJ64jDwKV5cpyAvJqLWCcnjxLr22zo8FC+B9t/GrtpOzSKEC2Gp
+YJq/b/St0jtkuwSe8BmWeWpZZEXUPW+v6XZnuXriHRVrPTaBfPeJh79TF6+YeE3n5W0CoSf5qVR
bveCxqHr+CFv7pLxVCSqC8fHq7dV7YxMdY1cH9Hwv1r0BXpL/S7M9alTuhesv6+/Jlie6HH3/nv1
iNmnu6lM9Jaep+YWggfGoevox8fZ3eJW6+6KuaO9s8L0NQLwiIC2SR1C91Sb4mxVmzRviHE52DmO
5knBCbsuoV4tpd/2MTenccipwGZhl7R/naw7tp0ifwxd826ZMCAgjNBNjsX+RCdPDDEkVZaQVknl
1VjS853aU1J8Ccmbg3O20iBQRj4JsmHXq83ol4cp1Ln5Z9ohxMkh5vRkWp6+eV7/8qYQ8RMRRju3
6xs2FAvKdYJ460xiXw7FBAyEDvy9PtH7YM3Ky3IQIjEYUFsLAvRPV9kUEF4KI+N9glNFS7EmzAOD
XmLBzOHYFH01FdRCNC28d6VG9plnkj6z55t6fDoan9q1Mi8atzuGq0ssvROj42CQgk1yltoHDbWG
wgo2LOTDew2fB6LXT0fy6YxAd0aL+hi4va9SYS4j+0iywvehx9O159msmzJ6Th5mZt1VDum8OO2Q
HBXaUoyWE+UeHeNnNwla2PZn3A9sDkYCUSFW4MmWU20zEGsqYl4Tb3SVGHjtY4ZVxPxRixknUTaR
qKRQqck/OR/uSkCkOzyTdoxVw5gmmz+iV06Z5P2kcm0CwOU08WlPMXKv/dkc2TpJ0aJRgbheb+9U
UfDO59RURpUaOx2EfDo4i+qc1+GYcx18fkNm5lI1GifEiwWzDbvcFCOu+yKwQ5hItOBSOwFUkYDz
DMh8I/lHgEFc5PXkmXnVmqXETY84Up0ZmYkXRkZ9CB7YMWQIxQDjoy4aV6gLMj/GoviJcHiuEKXS
YpZqCLKMoZnBt7jzWmN6kxiW9qkTQ3x3fSM96478xVDG6xWpGfi45s9WB0hHaAveq2eUwdRV4Boy
eUqI8Ssd86Oz7PcT40uJ++P9wvNIOhGSTIR9yoqPmhML2aJBK7J87E8NNlBMvd35w5nvfI4J2+Pr
txL4kpdQ/iXGXRiIiRGsd/gT699I1sHhJWFx9anIxgdDxaZHAMEKOM74VSNNaoFv3MIwnv39U2JN
/H2qgoBzWeFcgaM99slYAA5aAmb2IPGWP9roWg/D4FsVL8jtvYVuoV+8NvtbyDKO0y7vBtshR/wg
4WXB9zI1y/TGRARbxMc2Lz1ou9kupNpkBeAf1CwSQXSQHS1m0CnY6ConyAl5PjjWSW3pUU0W9L7O
8U4sVQ0th21d+FMMxqyH9N5+DKdhzLxRa0+mzr8eg5NxdF8m5RmxCSyG9KOvCE84UhLgTY78oas3
riPQskIPQetgwCI8w67W8ltX+MtDQsYuK6dqRkrjYYB0ryeEzqS8AJdLpHkE1kkUYMMciTyCYO+H
q5o4HzSsMaRdzs+hCaVBLI0VxkxyhCIbkp2WhB9Qi0lMgLVikTL/k2DWh3kwwB4tnyGmktSaOZ2i
UDr2HEYyr1yJTqvqOkBNEPNd81ZTbxb1evboi2GeISaq5XEQgdjD6z7n3hYdTif/UCrzH41GWNdW
GJzVLl4qDQgvq450xhzIhroOFupg5eZoxSHIkhIfTJCYn9oZ9qyVOX4Yr7lKlnJFKDRojsS3VbY/
1MI7bxhxgm23OyeSMpHIUEUq1QNy7Hnl3bPmknf1C3XtUd3D90uNqZgvXWIK3NGFZTwo2QIwT1hE
heJ5ZRXxyJA87rloy6DJpSP8j0wLA40MeAeKQKbDhL0EJ9Q0Hb5bcxD1iBDVhLhXsYv6dUE7ezYw
/xp7xAe0R2aXn+gvOndmQfHlait2kz1UX7lOpJKKdEmc/aGXLAyczIgGVT790rH0LBu2EH/yWnmW
VhSXBrBRDafr44RYaTgt00w/FckRlNaB6y4i/W32xhVfJU3NwzINUUB2ZLhzXQBwI03C6uASBQAb
fBnbLpSuq0QSRjLPLVZX9RcE/MivNY8UjxwbbOOcrHeGipmFKcQLkDXsZWjINirau0cDDrq6zrno
k4T8GeoM2hVWNprM5diJwBzNObU332dsFO5ALsKcRswpPol4Cx54o6xgLZ9hnu0M/zPsUvSlHUTR
xbSrPHHJcL9+aqHnvP/ETy9qe6XifBtY+Wpl4ZGw+CVVEwXfA5gNOuqidpyNqDnVLvBnfqJifPZS
/N2SJS4Vmf3FTVDKxocvk2DJeHLf0nhsM7MginzCjEdUamI8hPDMioWpLzj3p3IEoA4Q3rnmvw/3
E6/WvdBJEFQgVaUBWuN2MGvhWDWFZoy93WIXr3foW4GQ42qGLLdJ1GMw8lYvBGGZqko5tnDhvPep
5zaDyB87ZMmCxcgfsd0FKo+STDIewVzZNwW/9uhBVgCcA9w9Y2JlDrV4MengBHqtOnWuvRvPaRyu
fLtfidmPXh1sfQM1MoMnR+W5rdoqGfMDmN3w1KrrtMDvybAGwIKXHN1pEUNB6RsK5YY/j3kQSro8
brpm6RGkFCQ6yjDEfjM0O4HogLcsgGKYGPGjoPmqu4Dfj4mNWwNyMm6ZL3zogR3+c/c+6JyFzI0J
PU/LFmfHv2040+OgNUvjFB32d7/cbP4AYfA69QngJmlQhYKqri7z/hyrWSmyqvJUDiFtPhSgQhW+
9v4hsY8AdqSTvvm6zxKesZiHlmfsv5Hq58AundDvJ7/1+z4VOLLip2aqH6OzOV7vMpIju5eZCAMv
eveIyR7RhZoGqS+1ldM/PEzmvdzAk/L2tHkGBjyE90FFR6o3rgXzvdxlZs5h97UrlBxGngHImnRm
aMK1899dCeI/07z4hY3P6rZkI7EzQviqyrOWlZmigCVwlApsQzhfQ4Out7AM+AWm13fmfjAX2J7g
yfInnUmQ8jnfZUfHtpia+2Fop83ZpUIqnvqXju6S65/OP3ne2bqiKrmeoxAQzfHhvU6K3C9ljO2O
andRDGXufNlhrFvYtVpJvY2QK/2yMhxd3sFJNPXofnUao6CgadYgitRz9C4qOwhtcvZE9zPA2EmT
o8RadVrUvYYQAmzJliw2BE/XuZNDdbssxV5SDPxxG5zqvl3jjMTbNv6Iepf1X9sytOIR13xKQr3z
Kc8ErSDze34b1ze06PJMwo8D3lYKF6HRJkRR2g9Syu2lVE24AU+81pLDIu6BVmsPPurH+9al5q0G
I0uRwnIXuqbxLhFNCWjBitF0VjiiVmRyoCyqTkZplXkq75zM+bFQTqXYwE+8bDy95mdM0wBsjzTw
lB5loAXZxT5v1w/LqjgOVTcULyGs7E84v2cioJxjowKRSa4zR0BS0Sfn0iWtvBcvFbV5yRx/gfTX
VqggBH/9Bq4HoJIAhivgwJnPSQWHJa+wfpa+/f/RznqLLq4lWqzH20sazOwdujn/x9PQoCYfz6vj
4Nw/wsO2Sj+8iDmwQF444/gGtXRbHQ5HMNXAIied/Rk269eZ8gQ2+MgftDYQKukEQg9eVh2zs8VJ
clTlNn8V5wdcDDuWdgpfOHCUyG5ozxUl8au0Svwuhha1E4T7Vsg8Pf7hh7KKXe/+oz4iE+ePkb13
J6q9qbl8VcbMjcMxX27ey2NMvzWCyHe/Ec+m/cs78wjwu9gxPsf1ihNY7eXiepEZNu+31b9MuCIM
Y3s+ngq5a7/fuwhF8SW6N8Sra3PPAvfUf/X8L+qOzz/SDB+werSJNUBfN9kfQqqDZgegWOiuMpSe
dG+qtvIn38tslZeFsR2IRx4PwxRDeyTkyYbPFM/md0iAwUE627P7GAvDJJdrhhbaD1WsaF+Gz8mY
gx7TMcPEDKdeX4vjV5d3/L23lPCBC3y5BtHONC76sFCFNoFmWb1V2ZWdGJ6gsbkQEf0r6PMUh2AK
OyQ7mznWK23z932/pVn0IsgF0MB66OmdTVNI77zk2n+XajlmDnMDrer4CWwUF5/w4SQaPGNnGOr2
17LOYyNOD/E/FaJZWeGF7Csi1r3RPi8N0pizFMRFfkPtgW8CJZH3do4tNzC+5m2Dm9cBCZHn+t35
qDv5C4sB0ExuDNpI7rDO6eZWMUHvEGVA7MbhADVdVKguvdpiP2yU1LXSNdco4DQaLPVDo6CPQJoj
75dngbdx8yuGRhIE3aRh8wPSnwWmIUXbWQuUNzxuxo0H5hFzXkJk4Nh1koqPTFuYD+IS+c2fEHYo
XdwSh4aFxbZkcUleGb5Cf1MQjI96IrFJAtPpnjEF7j4bVQ/WzdzX65FnwnmAAwgQtULNXwQbUrXg
DyfeifsfmjoLEo4Fr6r7WfoNXtn4x+1Tifs+jHmPVbzbLhnnWnjYZV9gPdDD+H+DBHv/8GIigKrS
kYBDrPToeU8D06hIh9GrsQ0dKqzJYw1B65aa0JOnbZK6BT5KCAhDwUD0s/hqyWNHslMNM08+IGJl
nypPW/8EjQ4N/ElsimQ0tV+efuF9V1bSy76+v82vhkQA8siW3VYM2mnlKWrcToAVXobJyzjkyjGc
QMM1yrrTsC8Wbtp2Q5Qm3kpUYHJl3i6SINpxzH6/vZGcvwGrXrfY9QtpgRXu95N2TBxiW6LQaxi+
KgBJOSiRwO9IzZeFnaMip+QjSX/7gkyRi3gC25beQ+H1fIEM1LP9buLDnrTKfto5JzxNC3RdzVrE
WKKN7A0fx4cby4uhgSd5oZTZfcb5UgUsjm96Jepzjq5Pr4eskBYl2e/ubFlySnfNwUik5hbrPy0Y
HjfH0jksUfK8ZmcdFW435NiZGOUq+tmQwcD1p14PqnZj1aV5UM2Cm6u4zBWIrf9+hWmHinAreHSD
2W3p/jGV/DgOtLUXovog1d6l3vaZ0uxAc5f1B00jDHwCgmDxtpEj9iIH4IQzGNnJJqXYxkg/H0tq
tj3+rUTF+ctRqglh4pTfLrzuwS9cIhE+YYbbrSURjHdlYruUSdbocFk+aTXO5y5TLYf7KFLKGQ/g
20MH5j5AsNDVZ0uRCRsnC/7DiAVNKea8lKnKbacnnrrd3PPw92l6sSA7mPoQunV76PGC/61lwoYJ
JhqGfB5KOFklH5LLLUuW5GBoYFZUuhwSVKT+v2WUcyZNfqW0pVOympy+Dm/vm3CYwx84xDOYAlML
AWbzIiGZQZ1nNNdkJHuXK+OB7XWnW+328pGf/psEV4U2acE3yH/Fd1WB6kvCEZON0iYA/lI+NHi2
fGg9gRVs2kpWmsDrJXOHpbxfrz2VaV6CoIax5T86TiY0KZGUQ339lq3y3/ZLJUkhoOeaY6RMk6EN
byni6biIy4YngC4QOt8MmMTAPnEw8Q5tqd3li/jneAMnYjIu7TGDbEszPkWaoqvLXkEnpqBDax5q
dYov+3omX/a1ZcvcZjlq9iKaVe3bnsMWmcO76S7cJdmWg5j/UFkvBazVgP0uDgaKlibvhI2JQ9MY
OJc6J9C7QeoyF29LUOQAx9Q9usNvhOaRwkhW6hsM03lZVcKproIzDKg3HA4ZO8poqOuV1dh7/4Pb
c8o67lhRPE3BQO3KPNgE24WdVXFcwiRvpVaq5pqMqGZnywGotTj66sT4GVOTM+/0c0D0XEgAy2NE
n7cSazYWKl5znzyaEZV4AYlzIuayE4Iwh5vlDAsZny3VtUxDcZCxzyIdiSwddVqAgO7UzZB3wRmy
h98MYKbORqAcpn0dATyRbzwd/e4HQbArC+0aTMGUTQOQM/PzddwJ4a3PCghk43oocbcBu3CnGUJc
RMXwD/HsOH5UIiD9yVStiQBbuif1WwNZwd0wTNzesBEbR/eDns9++v2q1f3sFuDB1nnUUzrk7fu8
JhRrDSTLE5vE3wbHw8P5gr/yhM63B4a6+L04Mt00zably4UYK2r+q61Pm+ecADSZA8l8gUXgrDoj
V4rzh6rRvF3tzZwFvGuDB7IApTXfY0tP58dxsH7NYprLORjlT/M2ezzsZJVtKGpkbGyfmEeDc6d+
fmUfMrKVTT9fyh26Fjkno4UXhpm6TB/Z4yRr3702ms1sz6PoEqLXoASyCOR3KF6ZaKfaG45r/sJN
7kn6ijZY+kUcfbInXdL/Zj9sZ86BX5LtyvRfUYjIAHzxjTlNulXtIaK7CGW0xZNeqjwggpXi7s4Q
2Cmrk6XtnkEolQzE0zAydXYrXmx1La3HZthqBfIDcP11O/Rd/4DF6EAKkbBhcY0lTrfTFHFs2LWk
jfMgBCwjvs7NHb+cyIYGXo0RgOQY9DwNj6lDhUGiXtuvtjHRERKjeLyG41lH6vQuEpdOVGNp4cOE
MnsgtawfL0JQztJA7oLX19RA8XLAd4avEogTrVvm6p7iZpd/UMMgNs3UmwCqbqhohq0BELyGBBaa
Ww9V6wK5ti3NqyAiK2LV06tj4ggP0pMiGzLhVeOEbMbfcnGxNIf8V5z8CZRTje5jc+ZCAJtAagnS
zZxEM6aJMvYJN/I6N3cZqY49CCYRUDpvTUohm8y6JvwgMSuR/qBVJsQAPshkesycOzLeX5t2Ow9S
qw5jO4EoFf/va4JEMW0qA48gFfnPRSKNqMao0UHVzDNilrTrT9SGmWbQcOlMI6I6KJPeh3sduq8x
78x7e8XE7idM9v8wh4+RPnzDQ2BzbY7KRR+KJn4RM599R0/s2OMe9T00A/t9qh+Fcyjdj4nTTm3B
LqWrBgr2A/CnW9Sb15WOzjBTy9Btk9s26eI1d02D+bxRa4smHcAeTGo6QVs5o7hBQcHsj6f1XsQh
JG1VgTLvjZLWnn8lDTh8x5SMKG8i4kHVVDAoIZWxEPNeHZCNZZ4QtPJ/E3/p64EtT1fYWk76+R86
H+zllv+B5fHgUHm/DrPcnk4U97UVeZk1pxH7I2KCe42GTJImbZGBHrQcIUZgxOS6wm6ALPSG8qXV
t+mrz1PvFTNv5+kkwqH/9QBkztbVhw7RYL6iU7rddeaHUqkoUF+A+iOfLCxv+h0GV5WQvVSdXl91
TFwA3uY4db4C3TFBq5Yb/Zvq0EfC3B5UCCyC9KRs/CbSBYd0DcbtzVn24poZed2sjjCpjzRXiXTn
bm4MqzPQudKzPdx2dNI6ZPGXYM3+GdXkWV16N16N8UAgr9YXlxkt3bmkDhwZBb0c7r0eV8FfsRxW
+Zs3EnJK+QauZtaRO4pcgXYOw7WtXnmZ7YT3i98bHStUWreaiM/zx0jL2fz2oHBjqrWlP4+f46aD
4zHdqWyNbUuD9dG9mrmz3eAeq6DjBEkk0viPi90XrcYGsWzTZSQRzrDfunQXiEaz6QAJP4MG8o+J
WPUvvAvtCe2rT9qiwAoJ1hvrY2avecjCFN8VkZgUVAGrNVKsX8kRqwvJZAjncWHXhGFvul1o4Fnp
f4uDXs2UzqN0tK9969MdcPoWG65B2k6SEItPxi8FgEjshI6ciHez0CrvENVjzIw4RuD5qfw7hSSu
Pi0KoC/FxOO8yumqHj3dTxx5rCPnFU+fBYcKjsedGcsLh2aBqmiMVaC66jxs8USyl2QCC5HtNasu
yD7qgk93MW3rDW5MRdmLe0k34SrfwzYWcTMZokAOSjOqusHdS/0p8N+8t449g0Ki4ieyqpa40qKe
0HT2+ggcpCLMjf922pRx6ztQyv9x0bKCt62UDD3J5qSfgProMRXEDt2d/MwnwFC9U1//29jXQsq5
lPjCf77xPoKAPRqq02Es0q63pUO66COf7zmPRZyZ+yGvSQ2s+RLTjG8dapPN/sv7ts7gPMQ0KHQJ
oOydo6TX1njPMudTWC7vGaFdUIDM/M1UjVFcv5pcbfjLeZp4UuW4hqutOmnj8rDGMjAgjmF8GTww
ahzeLmfVYonLX6zzKbJAq7lA1+1tYWRnjff4UMyBcvVbfnOvlQpX0WHdUpJD6wzPOTVTZXhzGK31
j1zkZeE3bJMDQ5HMA19TSKq2eVRFZSq37/wTULdoCqH83WzfaIhcTaa6MefKPvKMUOCbza7uoFMc
3M0WorUvcTwrMo78daVoC3+yH4x3opcdiGM1OSpbpwE/5qqFAL7dUKHehVnjOD0NrzW9rKXzLpOF
ONqBHmZfqBsvq3P09w3WdIevK6c0uNzqsK1IALo9a31xudRKWM1gzAM8Av0DfQnzQnPMAXOSEKQA
4Haeey/Q4FMuxW/DCsASEVJB0jL+bM55nnL+6Ne0YX2wpkqODCa2SbpgUqz2LnYLx4D0qdk3sFF8
/46FRAf68FWZEs/0/ILjNsyebxjoQfoSdieM/q8nR19WRGzLiMsbiDPMtwCXi2Q16zoPzruv+7oE
YKr4qro/8s+u+qOW3MpVUGUvCJZ/F2If7DHCtgkXKn8J7so269lNRhUmExYwlswuUPy9wKHABh4V
M4rV7M+pI4r2FGItNOtT6EZybpluzNKLSJMl2sLUtt2kiqB7cFYGdl0MA0mGwJjKES28Al5FkHcq
0+BLQ9j/7M8v0p5614GeAivdTumJBwLslG+R30kpIIgEdpyI1Zox2EL0a7G8nJfD93u1xWlCBqEr
z8IgjqphwCEt8xaM1UGt+0qyblOxuo4STmEtEqPLK/qwJF6FNzjWwpFWm9490cxJXaMpByCBxyrq
4nJxdpKm7XCI5PuRvjTZ/PMEQmVmhgyDrufPUqy4EsLQrmsyyrFxaqfDZebeckT2/4ztgZtVh3vo
E2ivsB+Z6Iz7H9M2x3lsOWnHuXc04pyvACp234XxLFT1596WaqFeKjxNI/sKu5OY5BvUIen9YceT
q/N2sm9e2LkV22Fpjzr7/OXXYggdtQu7AhUNq90Hm4+hw3fcdqA5578JdmAGQJe/OTvxIsx+Y3Yi
AXakYS1FdNYr1GfrV0adQXoJVZX/E5pn6feY51Idonma1WSNSLs3Jj33ngar1aqxnjN3bhG1AGE2
Vptqah052VkoegI1pu30xJvhYubtZcoHB/uGyV4cUvgGRE+iHuXzXDWioKoYueSEQzg08oNNjPtE
fylfkNv2g4yQ2msQvQhCjEhBRvcYhzhZgpOWW/yALBqcGqK+Wjnxp+Ax37tjSrGsIPAB+8qyXQUe
Ogy+SkWdbuCvjzz3GnsEqBUEXXLvXXwzuB1WMGUSm7je81hXE3oDHh/qQxcamZB+vL3ZfH3w7/TM
IRI3jbYmrEPd0IBCLj2zwWkdDKqmFMTL6eCUHw1c/q/nR49NsINElesgGpflMR2S9Ed2O9t2Q43M
k42YO5360BBrElk83irwGrX91K8WY2bAwKBS0CQcXuVm1z9CtGaypul8TIyPvQwNRk/lQFdp9iv/
XjKCWOB/ejsBP0eF3JnVRzUhGThyu2f6PExBp1dJduRYYnQHf2fitWjAxChOL6C2pW+9v2R51h4T
xGTSkRbJFqgJ9/B8iVXPZDNDxxos4RyaLJTvLTVInIgpaLGFB6k4HG3ALmAuC5TGTer0p4zjwnkh
GK7nerSM1O6Wu5fQQhNe82tpJ0gf0Ml2YB/y+K0NTiJoLBUuuw5o7BN7zclaXLYZd5poZqUkRm8n
SmQ36qYyuR133ll4pzoPsD/PBUdwJykXZx2LWRCZRTfx/wUkysNp1F8WoDK/DdOtivlNSTFaoBMU
37/IENxm9upzhstGhsMXDU2vfrv4tUq+hpvYsGVOahissmXWpZ9CroYSJbHbogrq89i75tmPjDEA
G0t5JSqtbybaDWPus9odNA9jUpUb3FUUodXRDDmXifwu/7c15j+2v0Libyv6pqw4/6VpizC8QUmN
uBjp8ICb3QRca3FvgbwBf58Fq3A+w3dW8OeCQVBHvCQNMOvjPPGTrxKIv3e/K6ysHu18erR+Bchu
NhzXI2Y689g7bvruIhLyhcZ0px2kswDmlDOxcib2/NnG5CPgfZTR582hxSR65VZZ3SB0aNIt5oWB
7XnVyTDXnm1fwo5Hw4Q0X5IkTSNNPhQBYhwcIBGOQ38Vitb+jTijn1V7mihtstVxjR51/nze6aIY
32hVyGTbZCTac5LTJi/epW4gjM9YeFjR/2Hl2coBI1cRk6rcCSb/TIe7C/VnqEG1Ra1wJrz7drn2
SHU1/4OGZhrgapj2Zrzu45OLF+1GcvU1e/IeR6WJ4cy08X+TgVR88AjXkl2LBAj/VnPflq12iGgB
wgKuNjkyWsMpbajv8PbEItnHizIuJPnsulaGMsJOw+KJHOhrBoH3EMscnuaoGyMkj69PaUN9RUWE
j5x8t76YljkNC21SztaMgFjZj0vF/VwGxvvpzxI2zmWeDb1mUhUJm1BVxCTnQDdKjqf6Ajx9WUBb
RZUy/ZxguQMOTaCCECumt62DtfdsCqaltqQMU+S629yQP2DOd2h9DwozTs9WWQcR8r0ZJuINWBt5
J5YXOKCAm4hiWYEIAdthRs4m152yCm2t1EzKrbJGohS6mgp2U3dZfxdHDKrvekFz37vHzGha1TS5
UXE9/FH0s7RSPc/HcK8IVFqZCxD2+YFy+8PzDk5t4FBHbI04OyRotj6R3K7xR1tr5NHpoq4Lko46
phvgMFRZtf3irzyz0tHWn8RYsUx5UmnzhyGP4KKz8msVu9JOW1K8h6igeX65e393jvaZEA/2MYqy
fFIOYinTiXy3F0XLs+tsfEkE0mtRDOJe91ibO4udvF89SI43dNexCNS8+n7uOGi1rvTOaDHtKHmq
Yl9oAJSPpJgVPf9gA4dLC6xFm5UQSY8I3v1JStkTuYN6+mT03R2Po9Lhc40lbe5CQ07CaB1A8LRw
VBeFECjhw+RNxSwA6uQX3ftWDrHDwa6VqSzSQxo+ij+G7e9cU4vS23yi9dm3y+23MiDL2ueO12HY
ioWtx3z7whpmNQCC11K/jLu72xqquEDO1HwQ4u5gJpU4GOLHRwIvbcPYPnJ1OckOXo7lKQFZTg/4
wBrZiwNpKIN+tjqkd5CxpYFUqSCsL7y16KemN1fpSUh9x9Onzm3aOui5d9u197p7VGZzwNqPAEm7
XV6Er/LMJihrmfC6MnsMCVfn2LdVdVxjk/emjBJFvCMvSXtzFbL+QS6YwxZ7osW8fbTFYDhNkjH1
dQxK2F0dkHydSHhienju0yHh067g9nynpC5JG4F0IkE1LPGoSxoQgsonnv95I1V0VUXOb63jZICv
NZs/BBCv7IxbTnLX36iS42xO64+gpnn07Gloi494ciGwuXrEq7kSM91QD2HL8GJmgPnyZc+e5Ex+
PA4nww21Ay6eybV25lpw84tSQNEjUdYev3cKMkNFZ23h2Ld4hztvxQViqL3U44y/HtamEXKUyffX
0dfs0w0XDUrLV6QEgYKxnHPULIL5ZjUZQGLN1smO+ql8etbBIrIXO0YCe2+/boKG57yPeWnifarZ
OGAJdhln5Bp51PXzZkdVU/TDGNQvlVstNJIqOLzz8LTDcZVf9rj+wsPGE34DJsiub++b8Aq8m3eg
Nqizw2WIqBIHUGL9rhQkKbhCx9WcA3egS/7ktSqy8tpoxDRJE5gcZ5YWV9l6qvZl8imPgUtUQ6oX
uQpeGJMMxZaw78tcA94c+LG03UIOTC/Myn15Qw9nz0viEBq68WV/3tEoT9RlxiwDlkygCvMI16hU
9VxTAaRfUU3qO73QBIj9ZYt0rMGbhH6E18ZDTJnXsbhKQasig45+HPTkzrED+40JVdhAqo1SgeiF
UWShFvFiGd0YmJQH9rfLG6viO2SSQzyByv/picVIkUyqDOTX+qIej10KQreiED8nMtUQhHv3lt+j
0MUpvUSu5rfSpt1WRB2p9wy1bvOsJI9U+bHTT98abA5lFLEaQpRjpEy/wUg6AutYg+UTMXirLpAf
lqPoyMjPNvptQ1PLApUPt1YImwOsqlP2EbWfbDeD1d1SHNUV85E6xxcSH8M8rcBVPNwJp2JE+nmQ
iZdMLQi4c6ST1rHvbc3d420Mt7InHePlJ3y39426MB5pn+dJuNXF7YO2vcz1seoiVD3XxEcIbFB9
sZr4Hb+gvQnDPBzRr+hUnP8NuSyGJ/2uiHx6ThTx9zKDti5+Dbmh3gJmwj/s3Sk2dyXWX1XaHr2G
ByX/+NIrggxlRqyUP+LLwLQZzWYPJNOv3ohPqgjHTZXO/ckKha5DyM4b8Pz6fGUuecT7pzWYY+lM
zt11hyZ0aHIH7Cn/OXpINY0WpmCzTgivVkP0Ohyj3SeR4SWMruNEcbn7cvEGsJH5SvrXy6aVoq/C
YvPma54FQQlpVAvA/uE034lPgBkaMwLBrcmQvYBLKryWDP+uplPb3e1QZd6+fAFJDTAyuqFrljw1
lv7zLUzzC3/zC5NO7yeBQliAw9j2uWUGfJ76NGrrIGHK7Q7+mRiZbsoYawCzdWBvbXlVl9IavQmc
tZGfIS0WlVRNYdcNJ50ZWKNP6ni28JSF4TQarYwI2yRpnpkKiniP9fzN7gcKxY1E0WcbsXYkyrKX
j3aOIJoDubllY5YkQgJjEpH9yHk4RYVHOQRzA7sN954kj8e7UPqK9z+0oi4f9iTZgqVt0xd5Vcxt
KaX7wC94CTqzScUjK7zK7EOkSlblRG2bpOuge7n0YZlYktRey9qZMwz4otl+SDnh8/CbhOsCWZIa
r8lf14NDinmefKqh8NaYlHIhHijVCWcwBwMbL/lVhCeL52zgx5J+cJ20S/35Udt8GE+LcXAPgtVO
EGajZuF5IDOEl6t3OpIikKiiJknyLbyVfsjifUnCz5qhFSkOGJSsT48CyNMB5I+SYDgMkq8sF2db
hv/V5ChnUy4Yz0w05rK2+l+HKl/x8xn4ntmHgyHJg3PsCBzOSCmYcD8vima7SSiI9W6mtQ/xbWjO
YqdFu0+lN6gcf8YNaSI4tYsZGgH2Azwa2mD6nYV549kMuP+G9A7MrLqrUfzzG6G0ZEJZTCL5oSEr
Evpx2elgkGyrXOT7uwXCXy9QG4d/aq8TG+wFkQjXQe4UtiLLsWDIy+cDH7E6+fXWYhqLZMisoXdE
Z0hXDCixfUVyXuV5msbeEfhIHTuzVzZpj3WEA8+0abAlzzgNeGo/HqaOmnYTkl5YNq2XPqBO6rlr
9QooOOHhjmw21P2VDm539sMMjL9wLpNpc7hylRHCoV1Q5KHsDYMDe2zkhNOCpoOeXtxNtsVcz3nO
jHuO4XTzByQfQM5qfdwKEMOD+2sBG/D3teGf7l9MBOfownvRtKhSxEzCphERu4f7qOxRfi9PeY1P
lmZ+knwmbyBpwQE5W7oUBBMd/2gZpbPp3nUlw1Ps1wBRnxZO9wfc7LWI0HuoEOQZ7q3gwbPyalIX
fGyjTZWz/xDrZED/Z+CQqRCfqUJKmSxnhUSfmrjxG8o4aD8DgWbZ1A9rI6Rd3R7E7PSG9kwZGU2f
xUle8I38SximvNX73App9OESUOdbXQqIi9OYZ5Fcx9BFH2kOCdnoat+G4oCL8jt64RHoy/BI+TJw
5TpXxHsQodYT9osOWB5AReNc1kGUl3O1eDxxMAhONf6dW8x/1is2g/y8lHUIGcEj0NRNRMEzTa6P
94aa239Pg7VAFrwgj0y60lYURaELZbcAlg35ySVqVXGU+dkB9dEhwOHykJERWFwcv3C+GF7rDF0g
oY9SoODY+1ezGfluDhg+PfLY08CGzwCZDbD7BrpuE4bqtqmUld04TlLrDi1nJqS/fOBs7UzizK3G
aBLmjAbuJ7gQxzYnyK8cLVWYTI5+LOXpTE5BhTmYLwnCgB+lBo/27nrDo9XBa8/gsLYrcD6OATIu
gsGBaODOLoHY0ITrutvmYl7PzxcmICPdz7Aec3P+vgkNlRfXkgzxvMl8hZycWvLPEuIgw89Iyqo1
STZQPBPSCffPks82Db/bF+3bE2FrcI7GGLmbYtlIBSE1KYUfpptG1mm/JbGvhzTe6uzh78DL2I+g
+xc4SgrdIGSHAfydCA95wWfgJxRC8iq6CL8aYcRN5qkWElFWhcgJ2auB+ac1qvNiQMm7pEGLnr3s
KcFJCJCU2xwREK4QNckQnKADV+JA3lryEouPgFw76OVqAmh/64JzF4XlVW5mk8BJ9wRnIdm+zXY6
hN6jPeUk4Ts/K1yLJe5uUB43D5ap4bAi2A0tB70uB78h2FRQSqpkpiMTQCXoaFtIPTaanmEj6fgr
G0lGxCUsxG/KqVzT37MGBwOEhNk+q80ZZmbaiZbTeNTYU9Y3t9dcXuv2ebP51TC8mqkQQCo1a8Kc
WbSsigIiF//EUoa86NPbRybrmjUXxGcb2ZkTTZNlai8uzZvwJqqqccdEPTolBErUhsGp5p1woH9t
YgvH2mQ78IjzkGqGwMAVJDsLWwtv2IGYhyD+puiwosGXkthRxGfDRe3l4/U33WY40ebHzjt9AQ5Y
IBu5yLoQDjrtqSkf3cRrS9FCDWVgf65tvRCLnhO3OC2iOLmhIP/wvIaBDW/ybdydsAO0aTzweaSm
BNUKoQS5jkvlPpYD24u2S6zNR+hN5ibLd1ntNAxMMqMsZbWqsnw/9a0hzknqgAJ82Pes7CCzpI0C
s8ZwUbXUrrGUHY9Rinje59Dg4W3Co0Ip+4m3GxXn08nhlNWU6KVW3LrHbTDSWkdcxfK7MjtvXSDi
HY02Ib39ZAo7Am1ckgOsVjaYdsht2VxVNvjiLvmGEAsCw2BZl1OWs6+xxWhnK4QY+urMVEmCWChl
u//Gl9jvLU51XNXK4VtAFa8fwura/zb3BiRcAubYf7rlzMfJxE49a4nQOITaR+pNfZ0tlG8PimKe
b0X06fVsawIWTGddCQPgtHyOsCSTF2SEgeyYzyZujorcKKMd77UYo7BwkD9b8XX6oXIZlLrVuwFP
pQzjsu+cv4Jo9piGSID66ThXLHYD6YN5gA7raSkku8IQlQacr+VH1sYojWRTAku8RdaC/OLVbsy7
RTkrlWd6UiWFSSbvM6Wtg2lWGWhAj7Woa6C160UyVaNW+T2mCwmOKv29yI12dJsgucG0NYWSviQ0
WOZy40XBDQXvBnSB+3DMFVvpIPbNw5HVSnYDZGPASzecgNK953cq/ydP7Ti80/2Kp5L6lofzVW/d
hi/ce28AMFcp/Kd15qPj08yNJ/9/98g+9kbKZ3LGyY8a/xCEfHbWw+6JRVZLKu5BWJJgc0G7bSlE
X2ASC86PTPxv+thi2Skcva1JR08n6bK5BtwkAG8uKrFmEiORG+GPUKs2hhUrzjwU6wSOcaQFjmrm
Wv96qADsavbpdw5ihhmLO/1TM5iLW4WlJw2OYobMoMblMBS9keEfE9pcSVchokyCVbDSJX8EM0Fk
zl5PrucWj9t474dMi+rc5WucTNsoDuCgoSRMp+4VzE9jhALjaGOiT1EE9UYU9jhoBWi2RWDNpZ25
60fqj+U5MfO1ZrurPekMs8ZeL0lP+h20XgdXkz1hJewkbSWfVmBGDqGgwnyP2tBej/UWH9uovH2W
on8iatx2EuUpvyUfihCkvAwoH0hsv/6MrQSIjDyUw3Tsk018NgGHpVkUcn58SgvVGAzPQXzhZDA3
vQkoEl3oXm2/NFNmUrAWH2CRXjB7lypsxGB+Hs4N37l2WkkYf8RcJOPaGWMt3SnuVxZ4pdgRumIQ
janhcSKos6UhT0d6xOyX2qIJMQhh9BecN9+TtabwbA/L9ertMZuspuqr8OcQlaNDwKkHZzVkNBGD
jr6vn9IB+5EpoLtaMZPwHKqcgTOtky5Pn5NEyo5G+kO5qmVe/+U6I/i6m7xtKC1po3drF5ZpCIho
NtD7DvHV3fyLVGJahSR4ku/677u7Jy3nuJZ0GQosVWZdXSrsvKKZ+6e6Hzp6n+wQQ5kGNzifH4HY
QNnjJf3fIRxzcP+/DrQbulaNsYIt/AwPY9Aq3C7wJXXEfj3eOBcTiMVQs9k3oDQvDUjpZfJyZRzL
sw4C/iGNMMeJihIubE5NrEcsRRODNtA1gs8vprTKbq9uDes9EMlx6tpcMdOT3yxowrE2xDGOIpWW
09t9OjZQ8k6KxSie/biapD2TDXUlhWzYqI2vSVK4ZLAH/9wFKTuhn2HFPGq3kag//G50XLUs3izX
xnCoWJY3wOz8SBE3xpkfs1kKZl2zW1WeOYjjxb4FL2k3QC45RWsRsSRXbdNiUV+JV7VMkp9pVGgZ
L+lNorshSJyMTuwTsNv+WXsOR4RKbv04OBFmldHtzy5TO4QvtRSsQjcPBSoYGReftS1MTKjs5jBb
gEtk7xl1tDh75stCBKiBTGRMO5SIfjrClvnar3QVuiATz4CVz42kIAuQ1QUk5nxwjP/ZglossnQK
GgwK47mfLzvcCTTVBAYnnFYVvZKfDdpJAgfaQoJpZwAID4Mu6jsT77wy0A8KzmfjSlbLyoHEMbDY
lhMfqyc0q75ABHfWlwZvrCLyCUpaV4MQ97I1bSuaBWhXEcEA7idJk6fiXtLMYAfk5T4CICYYp/vo
jstGWaynqIRbwfeHVFOdBbRy5G7qrIFPIJnOaP/0szVgvy2c4eUBz0c4kGPoFvPWbKWcEocWMcnq
AL85exyEypdUhKNG7SS8IziDtJbQYv0VjV+uYY8bd2zxC6Ara6wA5sdl97k3HAHYrrRqXx/aja63
ihtHx7Yj0cLqUIEizbR24Zu0atgNW8UwFoWHxYuFpKR+WGATZ+4ZmdVArbhaAQDxs4KtG9fhFay6
CaarMLKdi7YuW5mXBHcPyTRpbipWmVibolPk3KHYJvZiC/HYfzzvgTa4fHF6XizczfthdDBwG4bD
JEe0bqNlrVKto4oFQrWQjEBFjNMcT+4o4WXi1gWcKXV/bW22c9PHRSFjuSP1i+DJ7pDtMBMcOmCQ
gD0+WKWfDFVkAb/rdI+ACT/kQkL+tofLzmOfoP++7ywc/O/RB2ZJoWakb5yo1ow1GFLNYNgaqF9g
Rppn2I1PHk7SJ1migZaRYfOhtVpD7I1D0pACyePyYRrZ10Qv/5Esbe4w94FGF1jNJ/gK5e2AuaG6
Ninr11T4u2pIZu6erInvJRaTLiRbryGOSQFGtUngye/F9XWnrPY6s1IOZftgJBucGxI7soahQ2PY
fMJJGgmUw7CSv+HJH1VGXO+/MYJ9V3RT7fEsFID4vlFD5tQAPX9rk7Sn3gKXej60h3BZsKx6C2cU
8nCscnPCT5Rduz/A6fcAZV7glRhemK1ZTOOOo+2ZHtO1F5Zm2i5QV0D1Zd61kMQrGBLxjXSOYi1h
1W/OCB5hTSuMCwbdFa1xIkNp5prq1QcnUqA61sVlkyBVn+DBnE04FSwoz0BhT+mNP52gy9Q9N/e3
dakTqUmDnQ16H00Jp+P40xcXeLubnWKMcHgr4K8ppJnVSCaJwxTzrjX7hVGVoMlerh1KByJV5oWV
Kub+M+I7rcA3F+fPi2LaS0oIDaNg03zRT08jKSyxjeTfGf5SgnZ7SYY4iH9eknsnwRIXzcokMDca
a5NYnW/5k51LbxJNE6nLrJLx3HIU3odJla2p4Aw5Z5HBFSmvLRIQEhZgZlWKw9PGmqBojMch243j
d1QyH1z2Lj6wh14adcTMZVkNWZv0mDtXA7gm943Y1qAjOx3BLOkrLh7F8Zx6gPu/l+S/PtHDZaL8
wbbjFJqcvJdFUrKfGWAZzr6wRHCHaNBQThm5hUCA6PqeIKCPuns5VfBcGWCPsmTHYdxf8YWndxR+
DPiX0LGCGaQVzJp69dJppZU4isP0NJ9282aVchkvf1n3NzcYmZZgRTQF83VABmh1F6cpRuI1o71m
l74SbgNQrFwidZSErjsJ03n9yaAzhtISGfbuyzfFSHKBybkKPZJeBeaBuLYcNBbOqf6c/Hq2YHKQ
zwTplZ3JMtQIpujLHIAo4nXVcZAe7AM0ZvePyG1Suw/WwUBthiYV/4cbyZGb/taEVFI1PTJRB4ag
zUZ8+olTAUD9TgbtgRE7zkKXHwYwlYbTNDYQP14dshGVIHVIJZdqbrnWJRRLSxcOEXIpoo/rY/RF
IoTxPh3J4xiILxOvSV4hTdWB314aFzF+SvEnartYe3sWf5ZjYSrqt7E/tfhh04TrwHFXje3MdBgc
9ViTvgWcRLSoiXh/FKhDG7xmPg7OqufZ8BtHlWo5r8gKrNIeVbjHnJpRMwisSXk+PDZs2RgxrQcF
NiTPJ84KPe/6IDPZ6noDdrq1mNCvXhq1r/fwQzus5/IYxLTrZeIsNnnx47kXFE7FzrZP02H0SglL
nL0tpt+N5T43T6vA6q026Y6qu4jrX+2lvSvF0QdC/VKjqV4zn7FDplI6Y0EPZe6RdTTSK4SKOPOo
4MHEUv/DUV10d7/PYP4CemU06CBNAbuEZx4fdncFA1UZHtNOppMzB5cWcEunAQ/xnggqXgpSMHzj
gVLn7HV1tOMnY/pwUFenUZRsRpd91fCteeuDB7apn3Fk/uFnKoIxf1dK5adaVmrI5G+cPW8xfIKg
FHFZNemI7fwXLYMklSWOGtXYuViXRQwFPjgde0H2q/1M+mb2ObrctBY055WH69vIGgI4OLHjYV2w
z0AFqVN1JDYO/yg4lhI3RHQjsQxqLVpH2/ot0dHzPyc+i3Ff0lOxdZeh+RWaJMiP0GgT7qy9c+XF
AHpgHDzwo0Qgems4X5XsPE91f7FKsx7QIWJBDdsRdElr8q4n0xChldQcFejdeEWaihi7P1u1sQ4Y
q2UNdN7qApoysepk6aTgf+bnaLScYtTGWcWx/5zgUn9Ae9nHYaDxS6E6eovZ9FoFmJ++TgCsbeZe
6yYnA7HkpusZArU7vT6ZUtP80ZejEV8meJnEqwiRZV+vtt5JaHNOKu1bcAnEr3ToeakJndOkO/lC
kWCrN2lxCM+8M32B+B10ODmVLFrfqizHDkPpWterLO3gW1jsWk3c0X2a+XXZrmD/cNVkOhJYIWKe
mwEg51/Dh0BND56WvPqRKmFZR0TwmK7ibOzomrRCPn47ON2QxbCNX60XqTQYjlML/pp4+VIuD7aE
rT7ICBC4Y1A7+KB2cLmOKECQQS8Se7d3vYmraYbK3nZSFHZ5xuplTJr5Y4tk6AqRFY1NypPRnhCn
T38urgXmzW4gc9k2Am3eJKoa656pFjFWqlcNcaE1T0WnSAV8/lxrfNH7VtCt/NJjUJns4OesRJzy
ZXjiG9tSYagj/L1jaEGQGK61wELwT3at9dTl3ymPl/NxBqkvQZ2C8qOuxHhaoDf5G5svC0vIpfmk
KZ4VwWtKBmVf9WPILaJyJSLmdoUxYFwBH3IL3Qo7DpNewA8t9hfPQz5kLAx55YMp1codg1kgOdsF
oImZ51gKygRonyHRU/El2vYNpzdFp0JKfeOgkDkdnecxRyzj6SisDIBNkTrWHego8H4J4oCs8Kea
dRYpgp6B7JCku8Z4Gyjq5vvgZfWeqDUFE8T4jXtv1emvefm6XLreE2qOOyTSfIufoamqZPhIT+1b
RIzNX4ezDem72PTGIVOhzt3SrOAI+cV0kb3F+PYpCsoysEwIznKs1O7CAu54XP54HIj3dyuGpRbM
hi6rfMLquUxZcF3o0ZJDkXAIvUPOEBrjAC1spBFE45CP7slU3dDGPx7m+yTmxQzzkCrhnklxC6/F
VVfpMN4trpyL/MCX4UzlTzVZbcgYrEGcUQV45g2ECW2TiwjvHmI5JNmbS9d5O0RbAxjdt/yQYkDs
WgwPixm7B9k/76RwH0jes/1Af3NCVhTB40PT4bZ+dEXODPwWq8h+D3+7xgb0POh6twuOhwVYoTp4
DCwqznBZAEcMABQdiwMxH9mdgLDbTXybw3VRl/Aps2qTc8vh8ATatN/UkhtraECUNu88ddkEgVmX
JBzEvTfdL3JyXaftsPy7lRSNNlaG2RiXeZOzu7PzYj58DZzWOTdgCyRz9G666C5+XjXRKogOPWpr
p2uty+AhyGOi61mK0Ht7fxUonELqX4jxL40TqjCem5GLtphbJKMMjAdeh4p96qfRTfs7KmShmSgI
U2E9cAqoOyCsIDAq57tfbTRFkYdnxLeTBwKwVmM3qEhiZCLQpWFZ4WAWOOX6PRAVEpIw7Xb0GPe3
Zlsf6dvRzMsQIr98prNEAOh0aKj2+cEOpHTFhPXVrRtAReoirMEAmzFCFQVb9wNCdeemN4nTdGBh
tyyqkfnf9U9k9aSvS7DbA2IJHD6otfcsTWveEfalVLyj6Am5n87+n/4dLXFciT+wLgTM6FpOouEH
ZAzQHUIs2omwP4ZSkXUx3UvqAU9TNN5xdjSnWMyWfxDz0P4tKjP3IIyJJ3oQfUpXU3r1syiU1fuM
9I9Mo4GGJnTYPxlujxdvoHtWUEhsR229A/1bMdK1JWprIcxCZ3VBJgR9V/yVksJ88LJXxoC4SvMh
XvLt6rY1VlAFPzvJyVj5bQ+ZJTACUuiE+HLol3E+efie+EQ0ILTTaDRS/ycgnSFODWuYztAsdSME
+Y4ciu4yTqRCsdOqWXz51HKCOCv2EoMF9grhcPjVSs95oSOkG5zckYAv+viPSb+oPjCZtCqvMSt3
dvCfiA3pE1OSpZ7S+knNW5DTmMR9JgBGs1VWSyYNkZcJrhXZlK4ng+nMI6E3IWZiQiVy997hcsHg
1jZ27/0x0tY35ciCpSbuCiFcYTyAhYdjiFvAitNNRiBzYlP9/NKjFH0ZQZXUvHNleA1CoOx3B9kx
vq73/0Knpa2RLQrsxsE7khzvPw5gKmn3qshpXJJbNh+T7gNoG6jsT3Spbjtr50sUTcdZFppXC1Xz
uLiDDvI3pzq6JEy4lip6tkv1f1nBqnTcItU+p1rDA8CEqIXM5VhZM85yitUwthaXR46aaXvWsPqU
jdW592HnXLRYkdkbg4/YDumEWKuRvIJe34z0w1vWiCHPKcrsKIhvSQwjS5+EoqkN2TdYSFxqKUYU
9W8g94RD9unFN/wGkl4JgmSu0sGQIrDrbiyv6CxwPW/O3QCL9OjngwWruP+sjNjS6F91DgLCnUHs
DnDq8bIE6wlinjeUrKld9g6AcJ3VKhBy4VhqhOa1arVVR4MgQ8EjkDqQ+2xLaibj+a+cQRK6LlZY
tQdska07Dd9QvcCTQMxq10VcyFoAwUb+P3lsUOgiTnAO4qH17ZCFXfrdUz2i/WT7ZlELtGiktsnu
gAWOs4ot9Qe2HyYXLeRdBBqAnXrtsr7i3ns9KHJVwfn8al793518nAX/NC0FkTgQ/M5iyFrCN8GT
CKGhGPv5ApzkrgIclXmFhAqrPpAXhUNFuPcGN8wIcpw4yKdcbXkF1yFTzC2/pLqS2yXVv4h70pUe
5s5dtMFtsI/rbNuGbvrje5/c/PJbi74AxJgDBShGpPLrS/wIDPMQGLJHSR0h4IPy/9jf+IKu15KQ
cFTQUwRbys9hSohhQEZmdd+ugT32vBYG3uu7NxGZvPivg0hDtL4msHZou8cWtoM+1AVTnDzzOMau
eruC/gEsp3vWzhl/hV+Ln9NsYVpuRS/tJyPcJSe13XriUKRFnM1QSmeBog9CsssQ3rOUcCuinUH5
jonNNztEPFCTp7OfN7wKOZixOKI9c/A+O8oqYMAzIqw71gSwdToFjXHMn43nil0sd4fsOwrDUal+
QXDkgvwuAp885ntE2GLH+7VFP3CeG2y7gwQZS+JMLrJRN0upEyE6zbM5PoJ2i+JV5RpyYk+bCLw2
pLUkvZefIwYQ8KQt8wdlN2p13lgaJwL1srl4cX2naRbq1LQ4TKQDysOy228apj5QZz0boOOXzTAs
3yYTqM+KjcF6Vv6umROOHhrShjWP6P0m/G8FOLOIrGLnuNEWClZjMYNgZCV+av7hmFectRlBzxxR
UQ5W9DSqEORiBhPFEgt9ELaPS8eCYJ511+MpsXlboUrzPK0/snuml/xlZUm9nKz7AWyNISFg6FXy
FA0N89zuFZH07L3xgB2gMaALs9mZO2KLkxCZSTxkuxzH9Afu//gyeqZMcFtt5jh4PGHFUCHfqSat
Xu3GMcMArrpobQ6HaYXX0Ey7/OOEiCnYiVbB7dMIF38EC/Tfaf3nNsTEn1qgEkHdsxFpgeeTOia7
Z/oYUdfDAojO4uf0WU+hmlAm81BCQlV+N9MyVa4xFhzkPM0BxSuWPGnddDMpmI3nOrjsiEzKJ8sm
sZJrBCdrB/0Xv1veHdx168yAJqShEfFoewJaxbwAkCT/7h0Wati90uO/dtJN0Uxo2ZyEiWWDVNa4
I2Bg0II964hGQgx3wDArb8vDF0c9UkPvFRVoCo8bXJznBYPcj7lCEw21vQxcOPt+ct05giR6JM+E
dWPngTLqL4xpioULlJAinovKrarMXi/zf1YYkkZn5zwKEolHcDJrXxYyntyr9q8t5JPDiUSImmK4
WNkZJzxhKW3c4Z6FrRd/+73hNQ3V4n6tyKqupDT7m5v6zaZsFfbqLNapQqzHJA3wAGg1cWhB2YyQ
8OgFj0dyYDg6/PIJzIkVUiSa4OX2upokWfIqrgTv0qO4RzTmPG1wRetO0LAJPcqqEgdoLhwBTKev
0Hv6AdEk+vlmWJgtSf/aRGnrF+uSBYQYv1YVklBdAQiaJr/HKoTqjV5uEmuwSEmRC5IcGQUGfZUO
Oi/IqjVnPuOM1UVkmiBjDbNO3GStK0S0Jv1Ew94ZVAcLIULa+DXhmtv0Xg4uwc0WRfiCyHAiFdJB
saAaIDHK+Yu8ibm0SPji1+4hp8heqt6VptswGCnqH8cZWjvzH4KIdsYNlZPk2rv0LgAiENdYhRqN
hvqmqMXb38+D24nn1yC6i7j5l9bkv2LWrHBZF5J9wScpFVtjozR87UqioAscGVez1L0SPBJQFPtX
Y3bDiMHqZq2S039s/y5KFZm53NxgMu38I7R8Lm4eAY9oFf1PU3XnRDdTF1q9hT7S9jOCDluV37TT
g9huS6xZHCuu4UAip/IGux83gGSBXaAKj4uVYrlF1fVE8buvSi6hv6856GRcWF7TGKGTIoYNZn/k
IDJw86TVvhdeywTfwDqIwmRkRm7yzJqwQAkma1mO2MAulFej0YBj5dRTBhPJSpVWA07RAsFoDnFq
4gTXdaNBc2fqKJo466l4GAohpIdteISkJyp8U8qzf30mlhAis2AVG9MP93aWKjuooGgYMV8HqV/p
zckZK+8AUtHQrpLi6vjbkfdnIjyYHY6awgTaa0MSRUhxeiVMb7O3++d3Yz7afyCJjJnMNdjiLO2N
5xHPu4MZ+D06nXirxbvKBSuBmKPw+IRzuKQC+Z9+gcTrIITN6Rlmd35LT9U+Cw5aMw2Gf8/kbofa
2lTI0TYscS1gy6IneADn6cxhUqK4JBbFsm1h2gkKyAar7UQWj/q/82p9dQRv5cgBlJ6DLS/GCpFi
pt2+4N90iD/VogL3zhB3leNBTrg8KiSQAPCpMi3OV8/1a7xGZikJkqFzYS4T3xqeViobVY78WpOe
NESKGjUCtiPjWksml6B/bM2JqyDKeeko6sP+f+pcLABjXfYzJRnQjoLh0ba5ZLdluy/N1M5fnsvw
hy+vYFrd8Nv1aSKeeqhfA7U1kyhjltU0L+mS/EmvH9O4vf+L+w6R8PVk7CMS9WFQu8uT7aIDBs66
i3E6HDx3tHhvxf8Jc2+DGjVTfQ4O0+cySq9SBEz3x4H8lpWBnMeGcv7I5UDTYXcxDMBib/+0TIz0
9PO/E/vvIMsfeNPhRJNtzS1wZcNmLFvKMwU5S3nKlAT0M6GJ6sqPiHAH9ik7aWbr8pMCkCbWXid0
aNZt0Ekqhj5FVfrFLp44Dev9Gq4NMzd2OWvfvt/UDpbOY7aOVH+VfdR2ZKldenHNnqZmgLY6kzMz
jYzUNJ/+VVti/+QMZ5l3izLaMdipVJJTDnV/amOyeyuCBnWD7RvyEPl82SRAhGl1b2rBVDlfwyjh
w0dQMo6BnO1lgGBvDWx7rOP87DTDZsmQKGiPW9n8GA++chCCDtIisD5AVANfmkrvWnbkZdKNdEhs
61qcXaRqzwR/3lWmKDHkAHbEvp5FDWKiTeyZZmZAx8R4qHzqvZbChQJfsjUG9lVhy98DaLw0GbjQ
7bihOoDXd44fUhjZtjzlHD4m7cX8HvZt5FgqSmpDOOOmfsiZEHLbDC1L+ffMt1PW7Nh8o71KD0ID
N02trItDhhL55qGymNhK7nhEwekfgF1RnLaPIkIRX31Rihgn8LZlSo7+D0hS91Hi8SH6rXuDRadF
N8YbmwRWwYORbbcEhMpITqWgVgMADvvmLYN4HBWlxv6Khpo1WSZKJxZ8HEzhOs+Tijcyf6VB0+5s
TptuwICLvw9rbafZpD+HUqTDggRb0hHm4iQBdmYQfkvlY48GhoNbvLj5trsu0IlQnzxRja9xgvT4
leXnZ7am8yI4dub9q+nZCjMbC/KKkpiYxRkFVAAB1eH7J0I8k7oeKONzW9o7VLB2fqmWW4P7u227
gylHNE86kQkC23fpw7tySan/+yQTpHr9OPuJc0+qILCUiAm0OLz9WgrCxx9UG2LdAWfVN+1sXPo/
I/hIZUxYpcOVx3Nfib9t2pMpAqONORMMZsXL/LIXLpzseOAJMjzAbu4alnnZu3lK5s7oyTmh7QFZ
B4WHXp4aJOP4vF3jyM83LBrdRWfV175QnkTpajgKiBMd/bv4a63KjvbQan7OeJxr1Zw781oNHVZ3
KOlfHGBWpl7DRrLyJk1dd6/TnJK7DOMRDr7T9gJFbrbDaQFKMauqoCx5aidB32yTFdsc81CBGfA6
tc3y0L+/1l5OKWYiUwaTIU8tP8ko7casexkKWAsBIomFCd6SqmTQogYSgVwtPDG7CGUr8qsfRY09
JGcFIQMrvhQjHR5+ZPa0sNeV+8sbZ18yYhTuZo2vZKS9NmeTs+RKE+eBzupyG68vZRKJVD8GodaZ
/JY/GtFwD+4GqsWBaMemykisJ9+ehcoAey/2vlI3549oFbj2LK8TxFSTAA9YtT1X+vUjP8sWFCna
6vI9enBweMfdLwRp62PGKE2bQ9ZyHou0r2lVnxKVK+tPsn8Psld5JlWK5doFDjaSmOZTeXKGyZL7
4XZrirMZV+DXxhhjP0mQ10cv07kb+FBfHqe4+cf7ZmonqvKUYJYxFDUfxjE4/A1jt+SPkBmx+sMx
nV/Hi4Tqa3BGdrOcqi0OADziuBfsOOOu2Xr/2pXIJcrqtLXGQjXUms8KZfGbc7uG9siIp3olpxZT
2WC18PIqEERVJdvgW5lU0QDUr1Sf4NxYZXbv08kR7T8mdvUOGynobQVzBqWpQ6T4UZ3VhZZRZQUG
lvZbKKnTB3gQkWZrWatwdgYdghdwXYdke2uYvnX+jr8iaPe+UvM9CWxxB2t5swkfWdRHvLsHBQv0
ONIK5s5a7Hc3qbzjG9ltMYBRr/TTjLBP2NXV+HoFbr3vvHtnZXr5VU1IAZ83Rmmi38o2WsZzYF5N
ROHHpkKkMcdV3xbLgWuzbRu7WE/SglxwzoNiokj1vN2zHbTZEqM7zAXjZtNkHwG2ULM7UCfBmweS
3APzZGqzD80483GdZT7MzvsB58bEY+jtifVnLxBbAEKdVuK96MSC9lctX7/6FOiKr3PtCxgmiVUP
31EvPlPi+NiwRUyr5AFAMujl6AgsgJOR0+30AUJ4f+gVsFUum8adW+iN7bhDDmHlvvP86nVDm7Sn
8Dc8MiSrGENtceYdHuSA5F7+rfJf0eO3/eDeVQJlGuwg53yQYRJyT/VEdBLQC4HNao1jzmKiTfuW
DjNW8igo5s/U9xsFAO+r1FpEyOK3DaYsLiLgRkOwXLJZ2qJ7WJFAAYhocu5LGrkljmDHpJxXo8U5
t0CsZFZCdXN7XJVJHKYxyS8hyikVYp0yDsVauUwXMcivG8agOrXnBod889TrlBrFQvtti5+GJ3fr
YygALCkuo3FpxQ1NWYQA67vG3m0Ibl+d4JjC/NCJVY/jVN9QvY4GsnJ0sEvCzhdV4zCwiKSiNug9
9rl3rcO9Gm2S9qVYGBRqdTlnfXvak5KycnIvIxfQo5Bdb/+tD3fMcYJwis7segvPEjIv6epKd/hK
VKKWvncOO2ZlOxRojZuGDdufczbaJJMBad64LUvVIH7KxMwI8jbhq2RWGM4e2QzpQ3VOQ9pgSjk5
sd5QYVXZ58kryziD63qM7Anb7SfqxgV1EiSOJdDwuGwIhDjcLB87GgFLCB7RGAz8GPmlKxkC3WiB
xTgzwNi2OgNLvmyxof35NId5KsS0yhrkrFNFUmvxZ1TIfjFDNjQFWnYomxeDIEKkMDCJHdWsTEFq
ZWw7HOaT8eDUqNUGhWMRG6LtwetqnENQtw4je8JpR5Hp27a+5qbDv6HYMquht9FKCRKp4jW9W8KC
20Y2qGVESXG0u/KGdAQoSOqlEI6JJPaaIdy4spDxWO8YVxNgewN0kJKGb+6hrPCHSYamEVxy8e+M
+MweENKK/GOmOgkqXw/sNaRjbFfThenfoJRXkJ3LtG4bMsyxuntz6pXtw7HOsFdwDEOiF9WPhU/a
mlZjNZ4f1C5IaGj32s5UI9GmzBeVLNOniBlrNlnQKfWW+oTk+A8UvUcdWpaJARgT0e7/86dkI3RF
e6cO++jygL51wXbgBQdwPVQVkQK7cfdvXwBPCu328ZT7oYgE04mzoZX1QDcg05Wzqf9DYTNH201k
Gsro9PwfqfiUppLl8x2oHdUFQ6oY2sWfNRCWylpTWEIZ7azUVtBd6Vh7STtzQHjfr/f8jqtRA9Zp
sAU4pDqrrfxqUQwKxKUUz/eziVvLlPpmHxPbYfhECPkGys7AvyCgA2E1Vx9XFs/W8qm0XVen/KAg
nZVDeMjNYD5zgaFZrZ8SJMn+A7Qqe16lpZ8hJhGhHT1mMR5fJPxvPbKLs6BUiPB1L6wIGkQ3z3LP
dPbwFcqkZG1LpCehFpt22nmfVCW/q7zHYqOw27hvimGbFcmmJCSXU5xCiQ/b2fb0Ib0+enw0f6i0
d1D4c5j7DhyjXYYUBT3Y5vWivpQiSnf5VRSvSrgHB0aKyYebCjN+Y2TNEdfBQIJ9LTYDog1zRGnt
xqf0RANB0HcYCh8uPIINzrRqIs7E8rIBAmmGFhAZtpNDpskSmzFsZ4wEqNVEEqAGLFkb0iAve+18
JbJLw2JePJ6subrvWToeAxzK6a8i2oeTC7EExLhHQ4s8UWzOfyTh5E31PZYDLfgCmafAJjtENydm
n8ghaSkHF0eEI+ukuj1HjdnWAtDM9iqUcX9NKN4aRyGiwZBi+opfQq1OGlwBVhsbXmhdu4fE1uvY
UBim+EpMi4xYzkbZx7sg+Q+22a+Mx9hr5NTc3vmCiud3wrBEU7ARS6xqb9BspUjEL5aQ8+JSm8W8
fAhAAy9uMLFK1ue0ZrjNEzddr4VdtBTL/zqQ3UbvOVDFYlc78J4JtoueHmavDd/L6J2ggE47AgrA
u3dj2BM73fhdcgCZw5AhEFD8CX2qBdwI3nGOnqvrWYwU1CP0t/Rw/AMoBBIuATPs7UWa7vvhdcF9
ReJHD7qdxlVKAI2On5yn4VjOALpvNatEy92/s/38dombZ4TqZbpz/K8aI7P74mmHUtyVMiW2TUBS
afbG6l1jG9uIdeynZOQsiI6nThvwOWpbSDi6DdtL9q9ZzBGLu4a7Br6/kXfMfdEHovXhyjRLR2DY
NEe9p4f7ixM0grFIesBWfdndut6Z4X2jLUf63PFqnHCQtIjRo0t4QLj5RBQHBCjHY0hxMpHj2nVs
9pT7I1RzZmJbWiBqYOKox8Y6hjsjsw3BHT+nNPu6WJqFqdh8vwidS+/vnTCakz5Lg/sGr89vvUug
8uVrx9kL4s60cAfg/apknW6cmVDV9tdBYQoWvMNROir6cVpcC+GYWFo1a6wXS2UGValGXdxpWchX
n4VfvuGNKxBTmKTTwp33A8cO7rViHh4AO2bKgniW59xMME0dMjzyX2rLHQ9kYDtKqCI6sNKjrABl
9ye6Tcz/2sOvetfcYsulRUCHqcumLjCKl9zvxIHSllcMGKzjEx28B209VHJ2UXs8moG5kk284wua
RuizkGVXqVOAt7hxzKdRQ+Wq4mG6ZVCFsmTXq1+kvRPidN6ab4mmH/+NhVUvsdtNqZWH1lzRexK3
Kxv07VHZkP+zh63N6z+q7jC2O8qamK+49eml6FR3Eje8G6sdwZ5lqOvwi9CJbis5R/Nc/M2EZEHX
MiJ4ndb6RwTW8ImIQM/XcWrsEwcd4IXNMpaBT506BP7oZdjz2kMATasJTs2ej5GkPEd5anHhO34T
kPsidP1q2Dn0k+ZjQDjXqJIjCb2QguRbRfYfighHdV019SoommJdEyEIf6Co2waq4aUMhs1H/IsJ
Mq3vLuhMZf6GijsPWqjm1gDhrSXNYgiww6UP2/AyztlVDcjc1CuLQpv4BCo9c0jdZYXT/afltxYj
+REHC/I7NZrk9fDiqcOZfgT2YKYuk8BNadN0flvQEoIvuqEKRpW+ujzMtWzZZJr062b1/YbrLSzl
UgoOQxRgpC7g9tSy33ljOFP+HBzy+7MBslodIbdDjV8MxKBHWMxonbTwsWTDGGVg/DDXigtB0cAJ
zYZdYRaSQZblFr+UH7NyL5CaIgFjSM8p/MQAApxtSXvctPe8T2vowrQJord1xDDZ21Rs0KOxnpPM
+KwiJb3NskHFyyjNVymuWdJNnvipheATI/D+/2uitqI7LzetO+jbVsnQ4LqltiP0NPTcnK2Np3Ti
C9+nH3xqYGdnhiHQBiJgZaXK/bnat2CBLqQkHcxyYAzNT1N4B+6oZ7Xy5pfpnfES85T/edxXwRSd
2ezeDSdRqaq/fGdWHBYnBrmeoJ8Z20PLayC6+z1HMVZILwG8z0Kgb1Qx48+KXAV8wvy0SIcGDyxF
htlqb3o3j9UIErnrR/hT9th1U4FYlg6z5LzNCMCJ3XsfuKNh3WUjDtittnirHrhcNG9NLAyQcKpH
uQ8fpQ/XdGNfsuZtEaVJ78rcRZyjnV4XwGq4jtZhmslFBNLQmQbrjGF0JuRKCMGLquylRtaHguaN
wXnKorZFLoy/63qhUAvxeDAnbS8CFDCBwX/MiqkwrwK3t1bj/CWbPz2moBkQntYzFJBGZZIx3hh/
IAAnXgIkggHQnD7eqIA+Pd2POwwQ1m5lf8PkTfMJV9rSpkMN5idLr87y1NqNMqFZHSeszAMvyhbZ
C2eOX4vZ43fc2LdkvFn0vsTkQW9IIkaBUT7BnNWlPLbS/Pfgr4GuRmCCg6RCvd1UnNRJH+FVbTi2
XLU/nrTW87BrMQt6KbICJsiermoOFJ5T0K0RHnq35Tgr32ILfgkN11ZMjOv7/oePpMQSaMVJi1//
t/gi5Xf2N/LrpvNE+hFx90GAwJsviaP4QothT/+PZ8FvQMAf6TibtTFCdnKYuGFfF0KNrQuN3g5a
2x6lHj3PHSeH8J175dVtqiPtPwfQlGlUBh71hIt6pPY7x57evJdPuyvMaN2iZq4roYjEocBPSt7V
F2TFi8Ke70CkRM3wiqxMaIE8cvCe7bMoXiZ9D8wXKWz2QU8yeWKpxtFbYkdx0Gp/QbJJ4xnHwS9K
vh8eX2yUIrum1r8rtHCw66zmrX37ifR3lZIQQIecVl6MASjd3TUA/EWKiO2tfc8PheEzoktForzj
bFgGrJekbAYlRVaXpStich7eudzuu/LbfBWqk4Yf4RUVrhuGYggZXP19MLStGoqgLe+h56gAr5On
Tpnlnu+9DnDA97s3612HuMwVVXPubVT9ZHek1zmy8Hjy90a5Ao3/hIB7RTOK+PWNEQRG5HOea+2u
Bxvyzu/ZMOkoqSYz3ispveeq7UZ/xEiNLDEjB3pSBZ0Rre4rExBK24sCeP3aaoFUoaiL0KygEqNO
w8Szj2qbayD4kiaRr+qsSlm6VOWwqdy1qPtqPmn9Z1qhThkBwItF+7R7Fvi+ut1/YTMdJ4uVrYcd
jeZKHfOmWoxLXWA7h/espubuweLU3bUJTWedrtRxtHaNBsFyM28+PuM9l4yrmtzIAaZj+VGgl0rS
jZJepK9vq/ULRX8P4+N4wCY+LSLNR0ii9oEekufUyTlg1oFMMfJQRf+L1GrrY3YRj3+oBJKkF34U
csadHqiSekUv9/kp1m++REwJActuBx28mns1pTfN3A9DJbFX648WhcLXE528fYSkon3KZ2Nryocm
74nNFcODD49nhid5ijpMxl6Q/8MC4zDS772Chthc7RBAR6a1XLde4Ad516Ywsre4D3FZMPFg7PR1
58Cd0IkujR5IiRqtgG245gmpFBOaBn9TeqWEUkjLhviH3uBVf4A3XI4emlm49ag1tm/3gIOQX8YR
QyHI/neoXuL5GmcD7FANL7WsVeIV7bc7JHKldxquBIAw/aeiBepaoityW2Ks78TY/pvTvc3YgU+/
uPyr8C0SiNpYgEaCCUOQuSYSGUEyIkw9rUZ4TtBp/S1ZaW4Ow0bxhs841icfx48Os3PqUM5qjsTY
CRypx0Bk0el00vdbAd8Gx60GliYNPM0NIadYJgVmorqBsn3olyG846vstbO2+Z/pA10OirKb4m9r
PPiffe73SybMgcS4lzrl99GuDWnjMZ02KZZdMD067zHcKlz4mAgyXonnKRYp0GihIGTwSII152Sb
ov3IHHbhzLq/10sxlsbW/49phQdJYpsC9prAxiybTUmjzjelk2maW6tPJ8tQrqCO6tajkqeg1oSB
ZIL73YqwbGCHv/jgYc66KVwmKY9h59vBrI0GSQsdotU6VP1bhdFIXkf9OXzCn+M+J6o6x7pUFcv2
kjx0gNgTWFjdh+p3P1AluFKFYbf+JzY3Qea5mhJTlE8Scg3vzi/fi0ze5FU6pm+1/zZv/6kLJpU0
a+h9eJ5wBJpoNR2w1TInUDvWYBVbwo1WSC/FDtnZl+JtR7Bs/ZARwobFt0VKe4L4nTu/dgWwxTtp
+0xUKyH94ntEdVeAINfl7P7cG5x5m8d53tRQzIEoMXinLVm7yY3TDyN1ghv63CW0z0WGryRF6ZTy
psjQF0QBtLoFnIgNQv1ZvJK4ks871itneRf1NfyWJqzKmcpeqbum2lcQzR4lr5a0Zqk4ayUNbd4m
Xn5mQV/KMCuCy5CYJEzJTM8zv0iPlBCHZ920eURute2lrqM9YMMf9KfAC7G3tqLjWw8baM1hhKla
tVpnmH0xNja9LehkE1ojINOKBuu5NU6pgaHBlVysgeJqhm+qkowjJbQelFugEafYqLzdbrnuRrka
CZRs9ovcR2KCPFANUwjzgOK5qwT6cRVmynKbNtDbEsj/6TiK8f4h1616rTnfXvHXSX/d2YPbCPcE
D24w3EPaVW+CfTZuVLDKlQqnpAC+YWlZt6uquyC3FhuBBWXoTrmubLTxbHUeapOyJVwhYv014MQT
yJmJu/D0GXYm+YQEIjtJNqXvAUspNLrBPrTgekzeDdeV7TwfAbqiSP35xUDrOvlAoLHO7r1a9KWq
7jw+FklQRbV1UZbgilMuKNMsgq0pM0aXmLx54No/mFUMd6fUeHadZUiwD+z4Qv/Blp4ztzn3sv+z
FmOM/qRDqN2KSYfFmi9uvDmWmlyQRDxHv9q5FxutabXQNuNPTWEQkGkv53F1Y0zpffLdNBUilsKU
URpq9xJhCGS47yGYaOtxNHkVB2ZNZsfneXPPVL97DvYaGTT0aPMzqAY5y5IQbAqoEo4AaEkW9D7b
s1ti+OxVa31RF+Cwv77RwyKE27Fc4xlpYb73fdTSGt1Q1eS0qrBwOUHB0K+ynS0kiiYQ77pMzV6i
995u3OVWVzYpio7VjuuOVdzrm6Y3vDMrRHLK8F7EzN5z6akOMRU949JaLUCAvZyy+l0OZiQHodTZ
VWFwWMSXDKtMPE/HWXt9/4+ttLEZshzR3Oh+LuYVH2WbKOPyVUCaxhh++Jw2uRWMlgbopdS2sHOx
gDoU7as1QKGGAg30qxlEfZxBUzaTaveCwWcmEmqunpoxofu7CRWp4COORsvHU3CSkP+IJsD8dzMX
okjBqiWC6Zndjc5QeuwiSrAg7WZ/MJ0lmqhWBXP/rrbvHLlP/sFcQqbze9xjWKrO+wxiRny4EMEC
TMhjznWA4VeOAVd3lns0sT6RQl1/9GqiPvMh+8NC+qKgHoyo0egTPRcIxGvTqybWItzxbRXWb6gX
EMiDTdI5hx6Miqaj2Dt3xcDlI596NHvYqRoQ1C5piGfDU4YLHR5ra2A87O9UxszzBSQd+JVirnNb
jkxYq0yvusn7X/zr9l+m6CBykk9ypO2RKBGMZyagYxvXmMANq6J4oa0G7c4q8iNNC136wLkwqtyc
Q+UzjryFa3ENOzyxg3uiHaeVeB1AkCcfRiKuLGjgW/19ZB2Z5vSToMg0fC7ZFgcYr7QQbBEOWQFA
OwsnydoA7g1f3/JREYMtIxI4XGeGq8ZhO2a+azB8//Dj975RZYmN0xKKGu5keeKXjdg9y1EU2mGH
xpiIdRNgT93LraX80KO+9HhdQGntOexdpo5gPP9FJGYriutEmo/HcZB1lrMx9GsBFHV3uPgTMnpV
hRNV2F6g0uK9H1/G6hM4tM/Nu9TQ01jjKLE262dGbO1FLWRcMLoeM1vHPB42MjNkXnf/jkTlpi4W
DVYtZAQOL6fcIAl+lMHtGWvBOUhayX7E3qdI+o/l+9em8lEGOtBqlog8NtxZlRdPCGzBE0CA78VW
XtXrZrMommX1uo+iJ1/edJ3gEFpY5/NHdM7yFdmTlmxyj330aH4uUtMLW0tbwdGUDrPZLlLTj7VR
d1TpPTidTBMcFlkjErhk1Y1/bDAr4Goerj6iyyOtvKwTkkTXX6UkFc406nM8z7n6hL1TeN7HLeNT
gKmQDc4MhcWmPbwIAImAf4wyIa44bhsfvuHqeYCjtMRk/yNvi1lwb2E1fYtF7x+9z4EwpG/YTvAl
7BUmbB64te3r52jEpR7L974eUi95QmI37dvEUuHefGvfIEZvz9UjcwhQdj956IkE+js8+UFzYWJ6
US1T9L7hiUnxmysnwqRFQxWuANyYvO/1tGWoUCvJWJ5XfLkuk/y5/glsR+JaGGratVbo2aum2fxh
xyx0nps8bYteaxyC+oqSRrdNd32ObmKn5f4r3QzlwhRejxMDbJpN5zP91pzjCngdaNFVl7jsr3Ca
LoVv6ReQ3hinolXu8udo9Eai+GHjCwJwMLp73X4O4WHVkaHGGPanwL4LJcVRfHK79CVOPFrqc0a2
uJZJHXbgYkKrfsYkOTKkMENPmmp6to95Qm/R0H+6NTWA/uJVytasEKY23EP50QkcGJTjJSdzX/Rn
HeSNy1CowE611T1ZOhkLzIaxOc0jWqsFfEUS+CkOol8Mn7hVu3lTzfaXp9LrkKC9otyd8XfCRaT/
iGL7gKkXcpjqpbUwT5S8BxvqISyXT9t59iWTvHD05hiELl2jrckm6sA09CDvIPzdr+p/Maa1TfvR
W8nIkxwsVWLbMCWk8Xzj7aaOCTFEF4nKgQBGVs4ulGUrCcHY1cntnJzVESfgfCa9KGIKU7pn65Tt
uZlraxfrQ+txqbtDJREJr+AGoMgKBQ+tybuqpHOVAxU/jhF/vu0ZxoH8RNzEggn4laiY2ru34ACz
ctM1at3rSD9YxG2KEqHdobtwwkbdIWAgBRiYVzoTdxZc+Yz+spFQ3ZZwageDBVnBQT3UO4kYS3WR
D25PtnX3bwKET+giBoKVozNG6db1nuFI85bVH5BnxFOuEjRpF2KNFLQfxua4226ndoW9dO2yz7vb
oF5Ay9f/GBU0BccbxbcJI9AUkyVQ1T2d7rnAzOw79656jzilHIC++E7Zyln9Kqz2GNt3muNcGtJi
c+C7wAG1HndzU8k1HUbQsR4A6Gx01kySNitlJBdRHY0Qvdb36xFnVloqiH7AFS5EM59y1FOfD+/O
kMcYuCztVcTHE+jPAlf4o3otDTjy+NtNkQtWjE0ZHkG9LIC3FYT83RiLybITVNo1/EBNAKHpMExs
8mXn027+cflnjkJdOM9Dt6EQ3ELOM08DG3WSBUULsGwlzvgaXWGGAGzHonOCtRQIwy5MrGs7nUlI
mj4+npo42uh+S+YNZ2tTj43icnPPpfnlHFnTIqPnhF8tk2r5DzKGMaTSqL+8OLnkWkSx5UwXOXzQ
WXwnChRSm4P6UDtq9ivFj3BNzQHd0mgkTVIDr/Ku1qNWzYqncVoxX3NsnQkcIRe6zz+XfdN2xfo2
M3RLxoeIWRMiNiogpM2YqNuOoS0ImKauuk4UsLWOYsCMHO7CPc1GVwD5xRnr5WLPs2Eakuy092lT
XdRg2BMZeqh3io1E1m5jbJbCyC7/4spMDx9JnXGi4KzFyITRUPK/PGDmKQmOGClOI/vkAOW4X0xR
O1VV8eaXPvhd7u3qLbh9by1u/V8ytCvBRbO4KfhFQY5xhpEvM6DuxDjYzjv6I0fFNFUNalCoYWlI
st/R3Jz6NRN1xP3A7DtTqtsy8onpQPXxvMoxdFLAJGaY6ab49PIs1+0XLCAyoNc6lILYXYk9M2XX
omUdJRisFpbI9yfhFKVyfFg8XwzkG+w/u4jYoG9FMgxQsboM4EpbjCRlfn4l1GhVDAffNPoy4XmA
icSqCsVMw70jfKy2405wJPjKjuMk/YQ3cFY7S+jHWPex3x/9zx3T4C0EoBCa8mR1xThdg2ceQ6bU
2ezHN4knGUZGSMfVJkYcddk/ovs1bBwAj9cLNwKDA0OPrBagWNm8uWnQpfqo5KZzk1rZkS0lj6B4
yhKOE55fXPuwqK666h1VwnPGjuz3pWViPsbk8Zm0kDGFd55mxokNaZC2awCL4krEEOKgpQtsEa5W
iwVhMIEOaNyOlMtIB+kQ8ly+CYW++1wCVfFD2j3286daxbNTXJhvSEh60MxyBnhmhlmRaxpGW9X0
yu6RODcGWDnWByyxkVFNVMxGo9PXmJX8mnCx2H+wliEBC0GaUVDEBy/XiVTVHG8/XFFMW0p1e+TB
oiy/edHUPj+MP4mFXLHdy9yuCNfS0LBjhGdZ7ZNztDBjiWj5GPJgp4gez6TRrnkjs9AoRqJeQgH9
0sdZ7XGRHUGRgBuYZ8ZlJo/KPVEBERSsfFmKe22c5XM1fVuhhBSc29Qv7SK26u99AiXLQ2AxF74H
mJM2mVP/YjQZja0mzDRGO1QJgiu+0+pmVuaR2iDYqeXH49k2+ycJ5AdFQPq+6yQ2eunkcgsL6dHs
cjQFDlgXXPOyEG06LFEw3ePVDs+fgWkdRKH9bokWWK6zNS7cTVcNQU5v8NU4TdCBMPhrBGvrkQcj
fjz4vPmrQdRkkWQa20vO4gY4RFBPtx+UpSprHDcMFUJ8NeCuK52tbDWTO0dIsGeEirmzk3TCA/K0
xck+FE8R5osinGH0u9GEUKAPoIH8YgxcFPJr0uPH1ieMzCrHf64q4vDxLrxUzKVsbqaq4QdzFPiG
1SgBHNf/iGYHlnYvwbRRwDYvi0xkXJG3zf2eRrCyZkn7td3Z8OJuw3FAa9tnK5Eb8T6zYeuHm2K7
RTrloIRO3wLhXSZp6o9aQpTDDnm1HK6nwZKKvvVfbPiL0hcXeSh8tVMzmMfr8Opw++Z2TWA4g1MN
DzBLlr9xu50eqCnpNY+L+c10IhdRpZhFJeUbkwnKh0LzrtLN+qsBafO66pLOuKm105i+zk5Iawb3
Gdwb532X5Su/bsXBR3szXlV6z7k3HDeY/PdJ4dWgq6QkoqKkttr7879HmUjhUkKAMfUW+JQoKoqQ
/tAIgHV/dwOE+v+TEmOq1/UjT7GyL8ViLxVrsy4g0zuUnDKJ8Qghf6OQAJ5CLaKt8DbLsEVqaOe2
l1gQAikdsVNf9Y01SFOZGMbi5oEqc4dJ1C4a8mDLU7VKl1QxZjB/zFX8Jjj4gC38WkTkrfC0TAJb
d8cid4tOpA/FopDeYJzKUI4liV/P5dknd7ZdOsqbauNV7Zu9RYD9jIWRnJaLmSDB9SkI6JUU9N4k
u0+o+pmmQRAhOGPX+UkgqQ0WcJedw1JZ6zK+VCD8R1bh/NXdYT0YVk9I/B5ILuiD6y610pvyu791
x8bQcxKfCDx++k6E3YvE46Q/9r5N8evr6ziE7jyNullhyNhzN5Y+XxzbY/UbUOIZous0NoI8Utp6
2VHxPeyuIu25q1R3GA1ZVNomCEZ6YGC/Ums1FnU3fbuwW/WoiUg/DqoPQ1JyPLdHC1ejwvNbyqRk
rOAIyeCNg6sSOBVn8XI0h64MHC5d8zY69w7ULnZUxtbBG8q+ya7fFkLoDakFcP+er695gy82o/WO
sNBBbqyaj2+CCwd42zOaUUVOrMJfIn6D5GXMUfHZfiax7TiV6cX5zjMGgR+Wa9VqKobt0o9Qn608
5VgvZJKWhS0m6SJr/LkBloDPcY+fEtuP4T7klSpSlGpL5MuPGbm+x1KcbkgY0DT5PLJcw4A5jUX3
CjqpI2+dC0QZz14u+mrdQFtUi6M6xH+m+p1GcZxrUJhkFqul5W11sSaTcR2tv+DgXorQQq+Sz2H+
HqrZlMlv+koSZ8LTNCK5Z76vT3/ynOO1jqOObwpF+C/lqdgtR326BTiE4VjvfNHvtUGXDQ5Tli56
468cNi5FrjBS0JIKd/6OoMDztJqcvX1039y57dh1jq1Hcrl79tNr+fL1BeQyurDx+olM+yEo1IBv
759FFV9ABEXjmVKwNazuVJ00PCXqiSTjiHamxTANRkwjflCVA2OCugv2gvvNI5OiNJpGcplFPrsL
cwZ8mRJMPjc2xhsHQ7GjlvLqrxMFnq5qsIk/acyFlvIV85FmMDJ1kWF3WoLLyTpvu1y6a+prVogS
YTlobwpfU0tJKeeqam6TvV3kWPp33JPjF5knObHkcFJNwREK2ku3+3rqFXL35BhQzd8f9qH/sw1u
nCqXvK0mu15aElsA66HhZ9tJk4CgJJKB4NmgI3V0hVbvKG73K2kziKG1C09uU2oc4fDhMqfXa7sl
wzeFkMPCIyt+rh38iXTH0pGYZdeZE+cg13GaRR9x+ddEgg/cCQbB1ryqlEjKmug/48k2ir4r5hsi
9lWXIUQh7KKT7pBF0WkbCXyIDlWSY55Cds2uP9dIxBEJ4MDZGNWlrIAmjHjZllv/kxXy+B+LCFJU
JaIaCtXF30RdI+rcxqlZO/ISL9LtdNc20NpwBh84sxrFeQTmDEwBe5znzBxy5Kd6x79SOwg35qWU
OXpChrz0cOc+kKwUpBHnPQKq+goTSRJnnd1GyD+ZvNCuCfs+Z1n6qaaC3OOTRY3aGzG1FEIspIB3
mnaaSwMk0kPCLI92VFSoRJnvtFWj4swsiFweL8vJFBTR0iagAfCZxXo9aiw+xeTgriuE0olFPxr4
PVDfp1CxXtcoes/zs4XIgOkWRoAwv5NuKQrfqfp7QR7JsiWEBUaP6cjJr/+CgKbBUJFfyS9meFxK
yKq0c/LgKsyZVtOpcNRUnPYjYnnV3ZuRssYTP9w5TseFlWVogUuz4R8/1Vnv3idpg5H45OIdyftH
jIl1xn1xiaUhgEy2q2gzD58eXu5qWs6DrMEdt9Sme+FgO0KBozrRr/y2OkUiMPCl6Lxi9fivdQlU
a0szxEPqxFq2cUQ0xRQGezNAvILA7RJtfuN1iv1OqRebb6nmM9WYfkp3KfbUAsca+ybnFZDBsXA/
7zliNq9ExoKs13DQ9MmZsAC0UGLIBwR+aIv2MvQ3EqDx1s2Kn2rIC0JBrkCEWghvZxt4owJRxG0B
koAj6hGOPuaSj/rO5vJld2zln386a/ttPh1SxVuqdmFG6lnxoq0nfsd8DYmBElL2FPCetmvBBs6C
K10dBFSwYYcbpj77kS9JSTh6NMq9KA+Er9FkiN46WE0iq56uUcd3rx+G/eYuRIeF4DKE352fXdN2
NRYRF17XxQXBrlUIAMLnGUVthuSHlG9krU4/3viBiER2ZeGEyWniOe/rIc1GUWKzA4AAWNvGyVFL
7wy4L1OD3OVNMHn/uELx3riJqYu46r/DgVWCMQWjmLc4GHO6mSRVQhRzJaEqgfmKvcZYYc1im5yb
28p5EWmdOu+eDGUjbLxDBC5nqj5Rwt6mEA0d2rP+QxPVmNsFRYOxQdw2KwimntW8C/KKWF5bEMmN
e67vlDSoHv1NsbXPiMLowC0r9Ix5677QotMuHlgdW3glhYeD6NFg6Tw+AoF3Qz+4Req610FPQr72
9kPrv1W06cNSRGvVnRcMnMIB3cHh/UaoOBYnTcUHd777wPn8MVdWwH+4yUULUmp0H6ht6iekrIDp
3VS8+413tbH0Ey85bFMqfEhVkbAnNZy5ctYEsdn84cY3E4hMu9NT+rChkKEndKwOwN5/LS8y1L6s
0NDGYxwEz4hFCwrXL2HbqU2egbzUiY2vt67RZiq8MhkthDWcTQ7P6dEUn0yR+QOENhWXHoCQuBgQ
WGfCCquavNZrXWQgkSnxJdqy1gwjEJjBW0yzFhSXT4Auvkg2DasoPqEx6+bwDgyrQUgmO7oNuGU4
/6puyMj5GEoBVJ2QJUAmfkU0RvZGJ/aff2aV+yRy6IQFjhsn7JujfBitMTKgG6TTmht+aNXo3I3u
FLjnk8OlDru0s7LhSO0t4vA8YrsBRwPrAv3yKJhCyV+CyS3vBkhRVruTQzEaHtZ1Kzc5J/psT++C
gg2WSKVK7FO+4YFUDYoHVkadUBC7YkOtYB5gZO0woAree3dda1J/KwlBmagWDqfPOcgiP3BkNpYx
iLR4+gFQwVt8H/2fuxlUC8iUsBPuD78uoGUGTa8p1js4jWU22wieoyt361zjlQUcw+gt5Noy0x/O
2oYChWQXliKlEujbCjuCvD+4eQeIXSUhdU/wzgjAEhAHIZUIOt/XdT9x2ZGRMXQKHq7FaySS0Mgg
uuAILFMUYFg8nlsTT04zdArQtQ2XkDL6fhz+2T7WzuxkJLv2xKO1SrMprj13BXzLU9HlvrqIrg05
RTIEKVGwhyrAuY6Po40nHDnwczjkePCKWFrFkHYbHvYi0g8rD9B7PFSafZa3vqCYZhMkmsnm1+K1
57WDuaBkxi8PlZ4rPLon0X8KRkT6F8Jj5pF5NUonVLqj9K+02mE2PvN6QG9I6ggGvpP/jNn9sxSy
N5eNWC74V49khi132ttAXyDpaiE32eChC0Fo/vTk+bWO0FfirGV0IzWl7N3RPIFDeAGcZiviGyJG
dReD7OVFwYr6hSj3ezcBgJSX6CJAw4MOrxpTDtTVZeaRLrTepKb3vUgwHr5GMoozc+YFIP3FUzC4
6kvTrCObznK7lxZNILkEMEZpFnzX4wMyNn+JJ292+OUOOoQaoPzqk2UjdrS/ZQ+XDIJhaTrAI6jr
fg186b/AQ3/rBn+7JMQTLcTiHa5vDVuAnBaU89Lb9TtLIcFfhVOAf8ItmtM2iT4P5lpRocWL6tI7
6/B0GLPtYkhhPH9Qg1PN8/kpvpJczpUEmUrfsZc4gUBFRNi5pPgKCB8Pl9Gpoi2urgMLr4LzTvyy
TOx33DGsDv3L6Ehtdi5RH6MMd1YORRqCzQPArx8hDqiHMuR9hbIevXJg9ny7XPx4Q0OghsTJG5ld
+e9Bg7551BdiWS5D/YSlFbavUaN2D6hQwc0NcWosx+26x/Meb7qfzs0fDAdLeDG494ul1MrNIxMr
zOQZw6wOikLaRUcEVqNW3U9Zz+ZrK1riMPXB5KkAManF2la2zL7dINpG1xZ3r6PrUDVgHtRtUqDI
rYFoiFP8tvjrCZ3vumYbymzSuM12BAyxV5VuvukhlKFQDjkAyhiacrzHW2pbcHF+ng6gzUl/h++N
4Pf0Ccl4/BCycJ7tkY3z3p6VJlqZyLieHo4KhebUjTZaUI1q4IlmrOVxhT8qHWGbrt6O7aI1dLKL
JP6Tfv8ssrK3zeAFsocuO35DWACSg4t/P5TaejZD4+wyZhg0dr7/OoG5V4JHqQfLodxPnAYTAfNx
53aCXmt5NMARXFecwqk3MEc+hdEO/awRj7mJqLygID9az6f1jQwtcXb4pGl66sXNt1lFzOH1FIDD
3e0Mu7hV4fx/TKmzA2xHKKXid+CWv9ixKDbATY5U7Yym7Wdcra3UFs8sRSdHPxJSiRe7OH1/vQX+
X+z+Tdgo2+ntja5MJ7ot5ZLA+sHj6Kn2RGrsqhgfyHA1eTifPbv/G88qG/izyQUtkT4jCvsrxnx8
Pd8+fKnLlNh5WCy12jH3SWc0lc3iVQZ14eUFCv631x6EDvepMVwePgw16V4jpB9xknguje20yyXT
sHtXfRItDXhXlnwxNzMJJclzZ5MyIFNukdnU0/tHBuZViNMwtWUT7peNgFy0dw/SbLMd63J0FAQk
3icAm/4qmtnJHHUEUBKyGy16O3DXY4vuDuvPZagjnt3XraP6wVa/sulvslwA9sW3lvlIyBLPBclW
Fa7gLzzs28oH8PePoYZ6yQsxCkbZkQy0kQMmsAIo+YfTwQT3bYjFXDmWLdprCxshVUjHKgARIYQZ
GwU18dmhUSm6WGQNRhPN+ngbFWIqgwRmTNLaCo+4u7SoLJmNSq9K9lJvHS4dV5IxV7W3k0Ulm+0n
YtWvkQCUiemuLkBppjsPWeHVWvPWMuzyNv/p93aJ5RWGQCfgcS5OzLrRWxUSJKbIyxVp/PM2U9E/
zc0Pt6tKOBOrhgSMThpcBkj5Oec6WYNyiYwhYgSdLUcrQuzmGZdpb1blLpSvJvqkFefDQyirFI7m
J+3mlWl6T1SAl+nlBNcPwOLo/W53mHgE0BQXBJ1PLfiNLPnXcdVLBblstxkqFeKxX8cPj6JVmYV2
4rb35jndRI3DDGlc/IivxyA3bY68EpsTq9l6d4reN9KqfIWf3yBNhqdfUCdcAUeY0pOc1G0aVBcl
VV96HapCeqhsTL2WGZu0D93aLlY/3IILJuJ5y2gkOyTYj8BY5K/DhDQn+M2WKgKp1pK3ztggVp/M
JKvQWGF9AmL/iy71yWRdNpYv9WkxE/ASm640gCO3PW8lKAE7Y9XatVncNMpX3QMFsxunnM9rhN6X
E/npEqBK/bNYsnWXSLq27/Q3vR3PtxuXv8pX+6D8v9L90k8uC1a+fFRsLPYlzFN2KizWGdXBvGW9
O5M3v8FNNDNKqIdg9NS0nvBaXwPG+w3HBR6g14Be4kPjooMTjDcdGv0qGJ7In9u/LVh2sr+pbYwj
T8jwu29af40zecUTDI75gpFREO5BF4CiuXcrPWKxvZHkHZxhtSAYD15wo5WIWn57LMMPg87TrJ9o
TKL6sVsOSEVkXqRoer2cnbuQWrvt0b5v+OmyjcoTDrNYisbCapuFEJNLbRnT0wAfPwNzQfAUk+od
/Ohdo8n7EYBKmLwEnEgYJoSNjTQ+kJ1RRbmMN0b+reT+5b19uQsChatffUqhYAKxza0KHUbwXONh
kmtogzh4nYvUbTtAT01ST3SzJE0w7wyE7ioPfXDtUf6gww4I7yM1E8L0AgoGXQ+h/Gz3ufdMZMXx
QhaiYCp7BraYf1y9lLYiqGNC/8ljIAzAaO/Vfet4AWB+Jx/FGLKyVAQFs6tyw60DuBbZSlKQFsn5
V9F3KS1Eh8hGZ8hwK9dFYYsMFLcnvHROFWLVv1bASqTUoXsMSENrN+/lsytbQvGbP/ofdIsHZgsU
6CFOjshCfxbpIwIklTGJRLL2qqs73LFtEPMtxQIre6mrBtlXYaAwAWHuweOqnyE5495iKSH8P0p+
/PijqkoRZRVh/CIMxxGNCwMrGHQ0MQIBRr5ZlYCjev2Dc6Xnu1ethJ/UYuJv86Om0HykS4/9uR/V
89vFnv+Nx6Uw7/B4ZcqbY6ftQXGCV4Hk7LSacPY/0l/NxRujbd8OetwH7UkpueTTa6UEZqJFLQsz
SrtK8M7rL8ibAQtqYONm9sQMZAnQE+Wz+FoeS7MVxQ4TvKbjZKWWeUfJ8MSWmW6lsH2HyDucpnkZ
5QZdIFBrXYJkq+iCLRNbw8iDvzZRPkF8Kj6hf0gONoc8JpgO5DoIRSXAj3fBuX6J+pmtvgCnU6Io
d2R8zgG5R7OJolVV5ZE4cb+K3bVXb55Di+DXNAG76L5N02TNC/ORDuVB0NI1Lx9wb11AEj44UFgS
SWSR6F7hc7yl0yBlhYeu9Koqu7x6m5CymfYvOrL5SSzG4vMjauq9W3ueQk2sS+oWtKMAnMazdHFM
VoIun5p00CDYH4F0uNs9oxd/GPkXvWgurzjlFY3Wen+GvUmCODEnQbV9/qisehI5yEy/TQOKzigz
g/FOmrX6RARNciIQzaXIKlOFdoA1II63FDah8ZYNImLdpFXKvresWz1Up5MKzKFEhvJYeQj+BPA2
IWjy6iowBDwo1wk+IpbyyqlRT/MrTh8NX+OUAq9JEpnQ+2AquFyTL0lshXiE0L1USqRdllIDfmWF
zP3Bpo4EwWn/VSBMi8dgs7rXGZA8AgY5drxLOyZAtys2KMYxw14JKx6yQUUQiL+vjmIjs1GT2JgT
bO/g/hQp9j2WBGM1wn3A85g+LGn6a1H+CfDCEzwEc82bmy9/iddSUHb5awBfSsEIAUzf1B3+NsE7
X1zXd+E/VS/5o/qfuTEJsI8I++3ImP8dCWixL6pnyxN3NGPDLcApRFHjad3UOljc8+ep7M198BdF
/nxGmzpKRanLolfBOpBPCLKGPsT2p+Hl2nBvlV3cXnGBigKV9uLFfSypzMT28JNntzsZUrioz6c3
fsS/QQ0yc36lqQoNycjCgTJFy46BGIapTH2KqgXqq8tmrG2Kc12ettE2axtJwkfFwNzq4kf4vb9G
X7LfsO2JPkNaoTmAr9XKKd43cj3ugPsIt7BsWoQ8lmJEnZ1Chz50Eivhbv3tIfT+Y4lutcuPVxaq
3z9oSrssza+UbLH4QhynWkyauyyPbPVR7UExqJfJWBRF7WUNami3L63PUQ6FuQw3U5+QqPHHUtUL
ybuzIXEyXRjyRh8OLhWasRgCqoRx3nuyQ1XlyI7x7WyfH4dBog9HNxKgxMsxLcsnd+Ut0cnoRyAh
X0VlJs+VgWmiTnTMWO73xUNTk+BRZbCoGMmtaqP+13q1gUv4LP2wH+Q5AQsj6FJoyDlfn2z5aFxt
A4OGWf3cH/ElLVBbFMSEzYxicuvS53cf0M9KQaic2uB0B3FIUzf45w1Cfco2uraGsurHtWgZRsfK
KjIvDg+6n6ojcTf7vM5mZz3o7WiORXqMw54Nd03DtBeMvQpgysURkQqWLjXE3CBY0KvCcfJKc/9m
RBqZoOqz8I4dEbDSGDCt8tcNgolSxGOvUjvufLGebYOoIDfFFr28hzM+a9mrjPwAdf+EWzUDsUtm
dR4IX6PATi3pTrxj6Cu0VWpC+WePzGCle9RXYFFxeWb4z2WmMnbM4TKG1fWlZDiIYYDzvIRhYAhg
NsBX9JJUgGw6IOoET+H7XjX0R+xeigmFoKxuSEEU9h8lLvpEHmX2IqVTyBW4DPoIgaWoDE6a2loz
MD+/BKi2x2Xqhn5yJ3nfMiqeivHytxcPvlrMEHVVoCAPoaE7NZtuZ8WZ7pwvPG1gnnXcwsjQQyKr
PDi1RzgiM06Vr0oMCMCOJw6AYZHxtayJnl+sFQWCll4zVAZPprPvcVCJGJrsVg+bxtOjftowaOTw
N+edJYvRnZOCrJ9ua4CZZS9ISoOAG9kYaMHj8/RLwfWEe+1YdzDYKsUK1LSrFKSO+IgVxkYqN60M
yljjs8O7oDy2ZjcezV0l5Ey4YXvJDRYtHkDRvpEYkqbhHkjF0INbiUl16nUEuj5f/kkY3WVQq3oZ
+KBn10e4ABHk2390qPtX6AbjJ9OavryffpvJ6QrjCvBn2rYGw+1eRQB6qIjj+jssJ0mEJtUF0UEv
/1Rn7GeUhwZat/+5lpPWFPRiExO3rVtjkyPNUB2hsSbD4A/WS8PVvrUQ/bTcXK55WK/htrAeLNHA
Mwn4HDvi809AK1OBfa69o/smLUOUOsLpSKIsynLZUY3psMmmCRburc7+TWVw558wSAdMDmtULkXw
mPvvhycxok0vISDNde7j/Wko9O1Uxu3nMX7UqcGLF+7UO83a+GLYUTrpROB9IqYVlhKgD241Xiig
My3rneOfnneKWwEjunUtPcRse4OsNOcDayGb5WAnov9G4fyf8vUL7MUs7VlxFjHjRwlXG4u9krO0
WL+NAA20SUNpSsVVLcKnHoy4yKc8gh3ZUXDdO+LrxSyqdIb6ocM1onFPabfAXfUo4OLORZ4AaaSm
4S923vc64MYSbk8mPUPBbyIGn8movlzoxTkEv9x9Jb1ahK35FuwL3VmmumkefxZohdZd6FSj+vY3
w0Xg26/a+TYlxbWPV8ozoafzyq97phlwJJZTbyspPoUDbUPHgExGlFT23rWg6Gq2zSd//s8RGwiv
lXpTQQylCioo83tmsI702hHrrpGP2Sj7LIsfXeFgXA7KY/eOaxhrdiH/u/Y3/htTIFlWJx4/3sjM
1/+hbMDqvz0muUSk4m+Q/riDdC/pDYUWp7VIQ4iArIlnMpW9XNuKi/oyeYKKaSDE3d6ii1DTaPBw
/cj7Gc3wd6gxIqhNZIsaetFN8BVfVnCg+sSE4F1Rq94XPUtTyHm8jSLkRgSevbCVwJDgDpsjsFNr
q7SWIN4OehfrfIQa6VSIOI9dTsReLHcKhni8RiY99/J9eLqh9iMSNAlCLNvFFSkiVDXgKqxaEEuN
rvCmnYz80BEyd4AM5ezNQAxomgLZPRKWXQmptVTV5sQZAv7jbcQeitv8bNGE6XfEnOn+QLQDXFh5
LvXDlMDlNmJTCGb8KwlgL+A9/3tP4TiUHdSFP/yE0PRiZFmhJ9Hor0Hge3tu0eFLzKqjiA8wF7kE
fgp+vXbPvegGWJxNR/LJCuVSgRrtVN6vFZ25O0ovf/Z9UJLDIU8/EaqjuhzqZicbdYkgvv57zT2Q
ASgLlMt6uNPCWsKNxI2uW87KgnV6BB2XB5C9CNSNQHm8jxXAkD0xJc4pR9llqu+ZmF9vQJyYrcWy
huoq863lYtsRdtBCFrGZ9LH4n9RhhcJJQDQ+h0/yQoKSE610ZTFJJtBGCVDVg1kiK6sQDFiyVs5I
SDKXNuRuCUMlCb+SAyw2lzJ3gQHVg2/g3ftBsYv8O0aY6Uz2yABEJjLwuk+Audl/VwLr4cCbmjiQ
F/ulgLlg2BBwi91I36ywVCKynIQu6FHbCJ8z40e+vY9gV4P2lF74WHYMajxhwqDtHrCl06xuKnQj
816k+g57v0NQDW1HEQCMrHK55bi3Tl9krmbRavkItYOdpkDjNPGvChxQr10h5RLvWkyjbG1o5Q42
et688IF7Qqug0Pz1hozHVm6xppj29ged1sNXcE95fxd92XEumHjwnS0qj4/bS5YQuYfe+hE2+TcT
wlHqkkt/Qp9npndhmfYs4unh/+9G9GO7yYSJNn8vgKGPk4wB13ii8In7xjTCiUeypcuehVgGlMDb
If3YmhPosM4tASfE0fZOJRcXeNfubFzl+S1c1x95r/kJEqxWdVxCSA9DE9EDT4FO+Zf/xHIbIlV9
J7AmoRHc7I6Pa8kk5tXI2FxtBbE/A6ZQWm4XDm1h+ooyA6of+ZwG/F0nlkIsr5eC4GBAOJNkqqUS
UvuFBcds9mCVcJAvtB7HdVdsiFG7xgX3MWrL2P82hUTBr7fEY9cpJONKUvG6fbuwmcpjwm3bAUPt
JJwapsc5Cbu13acD+hqPa6iRRwkr5FpdeAaK7xpLsSWlF3l0zbOpL5SZYTEIo+Hhgi0g8aezwfWn
QEKv69Jiuoh/Fv2fdFXIf2Il/gF7MPPhG2U6ubBogKxNAjoP6m0y2WVkIfaYAFA35H/bIR7dBx1h
2Yyeck8FfEfwIVMHgLvXJGX+/zg1AGxo0SAjxNif1aKvvFiQ35i5QnEM+9e1zQ6kiUujo1kLsCF8
iSYDCPu3Jc/KCCnU4xOrn9cpZUWGFLMXRP2r8zrvf/5qnpQ7kc9vCS9CmX1/ZltZ31j5piVsRaqT
6Q9njjHmpkLoBfMvfFfej6R5TfZ+b2pLCNYfqk0p04FgvRKOIDZH4X9QbNXdI8u6IU5DSWQEAWyn
vwn3c1l1sa/1xna/BjL/9MMzi0JV85nltQfFfhnVVyV3V4yVivlKa2/zClw/nI9TFUeRr5oooJXl
kV2EXA07J2kTyQQxkS/CyyARktuP0g1sYN36APISNeBU/Q+Bfb0Y3mP2stqgivVyQHUa6NxGhiXK
HcsHS+jbSrbQAdb2cvMEywza1Op9QYDpBe8e14vui/5HpoVS5l0Y/vwxx0+4D/grWdJFcqaoF0UU
N0K//zMsFxhPZu/PvEvH/qngD5KsE4LPNWdPIu8uLltpJefP832pPGjSS+h0+J9PZ/7YXktfkIYB
OvYHTJlkGsRVF2k4oPnpf9fWOfmuJ2gxIRKG5ElGpbnktTrdt17wN0v8ICIWMJ+m3P1Nq2cydp9I
i4VSIIOBUweENXfcbnKEg/W+lKa79b7Ok8B7B3b7AR1orX/bUS+AHWkot5lmhnAU6b51xdI9WQ1Y
3G881jLeeWb7m4lVmTGcNKHjlm4zaIbDlaI8ti2HKKOZQ6y82RDmOquOmHF5pCjeIcHrr85GjmM/
jz9LWMHHR7AfkDyyV2fXN9i/OjhasoUdTc1L1J0nRfmKaJD6Wo5dDaYGU3CqkvzHHiB9+QfVIWvL
LYQG+TmAv9RKYFnzVl9qQHvpEWQxKhHtGkq70U7NEdq6eYZJYRBNn3oDfrikwqoJpwbJp3R/YUlp
OMP6QKiDuZqG3T/gsmzgPX3WAfbuDJ3u4T2rhts4RrHYvuBYmsxABCPvYqhLJoA397JRmzrmr4RZ
QTxo5fy7Fn7529yFmp5WxuGlSShRSCxKK2AYdrah0L6bh+jYvmI1kqjevJ+7yfhOnke7bNqLiz64
VHwzdc08shPEXBD8J8MViB3+tpJxrpPpB6yC5H006c8cZHsTeG03QQKU+ChX5bxLeY/5jIAGXYPj
gCuQUPuBpKLOuxYmksslKuxRtUiSkgpYzIYXQPKc+dBGkdXvkvcRIpYX2kFnWjDrVuDxRMYz4AzH
QotiAtoNl6qyxY4pjdw9NWjvStk95BZgievH9zs9bvx7C+/dJjWevkQlMOygWuVIfmaC3S90z30s
L0tMhCUKMOByBX5K7C0eA9ccMGyJCRGqPUGzbdlg6ZznHYH3tDgYGVPFsjfS0e1g/O0FGs/mgYYA
EV1Vq8VbJQ1Jav4D/SYXJh9202p4EcAGZLmYVCjzLOUM+Ij2wOpF01PGSg6jpSelZ+ZtLMiVseP8
RwIUDQfBvrqhMExDhrfgJWCwB0nXTq8D7EVpet0wFGMjdj43aU9z0pshNKMFFBp41VgPifvAup7G
RhwMWoIS1SxkjSlj82atqgChOIo2yAtYRd1KclnDzCPA43gndzHNHpH62i2yU8leGPAlW1fQaHD/
50ZBvB45XF7+9c+ldIJgc9C/ZTS+EkNAzRyQYQxLN1VCDX9CQsqw2c24WJUTwa7pYEfPLRxdCOm9
dRRCrXQr71qbouusJTtWswrYQlm71RdZ23VCV1uYnzsX8rJGk2aofRiONzE2iLVP2I7r1xvmiokD
dfDRx5UPxz+nthqLSp3Lh1iVGOacM2u2y4qjAASXNewqPwrY0EJj9CPWpla83Reemp2nncYgXStp
QBsEUHT+sGJRFs0m5AyRQyASezcB+VHRdT/bqipAZN18vtGua4cF5g1A95kXA9XYX3FHZWVRxGrB
SxAWudLhmA8805jhBBLyPGA54nbCe3UobJxYAKltPwyBqAzCFYs4itbkW7Zl+fo+FiIGbvaAv4d+
AyzaEZLsqWwb1+pNIid5JEMIn05hTI5EseXYR5tzlUeiZyGr2MPGwNghMzJ9+krHus+QnmRx/hJB
+TAnhWVKyOzghtVnwQrpoOsBFl3xtyf3OoUSEeGoidWAiPP7/NVaCmTw6NwLpNRj9Q52S0+nU6bj
6GsKAwB0dKuiPFQc0V/ZTHqweDSGqspYOfhJmBpsCZsJB8FI564Y/ot+wNOroXizrJx7xG4V1xBO
aylrLpz8+2XBKjdZYOkqK1LZssWajjAAN6r00M+uyHeFSqmUVDWHrwPUwNQr29BoAlc1gM17XOwJ
VoAYa1Jmg0Js8NHupMfwdcqLyUgyq+FdFuNLX9wXm619XxCw8aeqF43k39Sd29zYokeAVa/BNw7N
ObNI7mREZu2LV80dSeskcNMHI0BvyTktxQj0FRApLti2kct7ELy6C12fXy8koerwfb30bDR76VRo
05s/UF+rZRP2L3G5DDVR0nJjZJkpUVNyTrGfxKYqwP3xOIqzYHiyOYkOU8sb09oTWJhn/LVBZ4qc
OfrmdnDzYha9TTvRsMKzupHp+i2QPN0rAFRVe9a6ZlYtvT9qcDYOMxzyxQPmi525L0Sz/C64vovB
pAtSh+E1IJeHQ5DjpvwTbn/GJiEYHJpO5Vcuy0AQH5sJ9mWqfiHRW4VUYdPh7dRCx3E16eqltzgU
Ngx6/0eV+ppPqaNsubpl1cNs9cinui9mlGTMmkFz2RaRTchSf/E2kbIwAGBLaCU3n/aA+nc5XXcT
Vle98eq0ZlyHRtuHgXD+93ps7QCrGOQKzVRM1EOOsoRE9M+4bqvWYjrASpmu9+e6vhUP4F3ovT1T
t2s9bMZ4iqVgD64NCeOIk+VEuAJoA6yZlZUl2m7M9+WEJpVxhKVJq1YyJXdYTBLe1WPtANa13uu/
swLipMsrhSKqJpJ4wxWM0wE2xmK7s67egi8LeAzmdVC7dYMfOUoP4/CZCTKAKwVWv92i6XGS4o1c
JpEap8imIsc3hH1sO70ptyw4MfYnclqNu2fcZdqu5N/wY8uTCDI6b+fRHZG8f8xYAYU/8MEkWpu4
Ud85q2Nx+wuONF5ICMo8hJa5IsX3ZP4wSzfq8LH1VDP/vSHbw5U1XKQRXsLuROTMj92kBOc8ksGf
UyRwtBYxokdNRUqVjJOGnymAsCUdfnuoM+34AqQ9r/UM/+6B0Kf3Rc+lmLVnSLtRp8iZqZWBFx1s
dB4bsbHyyGnOelnJin+L0YN4TjgxEw7IMNE8RR5LqHAJ9l+BK6WKilQoWZjs9D2zqg8fgnawjbSm
8hSgWE1R5cnLUt7FXydXv+DezJBC8fsEoxyYJhbWSkxYnhFMREKzI+X0KenQMD5pVfxSLKIPXyV7
4S2PZPE4IbvQVtrotpaKpOyxiM/ITuCZ3g9xaUq/7t1E7r1oIzaXxmS7880jx4Rusnb3c7j09XQi
Nn61jnkhNSUdM5MJDZrIiNaA5iEZEobhpHFg1gk1gJ/IwCn51iX1m7Veo/bJBpxiro67S1lmMpyH
D+yHnuZElYl09NHXR4Wx1MmhRfE4kOycQ2uRMyHZojOJiFEc3uBQLN+saDQ8Rjyv77TosinNAH1p
KPKhzHfaaMxHl3j8DaGQBFh4iasoSVarqC9JNymPI+1Tp+nlO8niHksRbWejA+rhBlKDgNbvT5aJ
p5zmTuc7LM9ctDoh7ws7N/1176sRjeoaieQ/zCdtR7HXyp1JQ+ehjMvxX51sSOFVweQRDQUB+BKC
YU8ACxf3vf66OzkXEDu1Wk93/f4Ho3w0hUsl4kkHVp2/13Sxq58HIcdYRTsEZKn74y/cipbvJ4AX
RTo07TWXhH96wvj8xfErFUOK9bGBFce/CXV0x/4n+qZ1UUQ8ibc6rtNFlvnjH5ak9R2BIiSp2jKL
q53UfMjFqxsIlgQ9Y5KH5zhm0EVcWq0mFCFALT8M4BEARRTPstQmlAOJWYLVeYhdy3sAmiI4DHxc
i5/LRprq7JoGqZuPIlaME+n9VXV+5P77P+8qS6gkI2kM9BVy5psfKZqqLR8G596gNESpn669YS4R
5aWXHNS6dw/d2G41nj0ZH4bKRpqve8ZMLRDs/mHLXVlwrp2GugfnF7TfjcwWV3leQ4GQMcfnqL73
UTn1AN+lbDjHU08ymuRHqgtBmdutJKzwlom2IF7HlvmQhbloT0JyojdJMaHNpKw0JD8HIxe7ThK/
T44QXzux1x40lv9v6pal1326eWD18gYO/e4MH+WCaeWo7Y5T/F+lYU3GZePKYAudoU65sU24+zqQ
1073abSqP6P5mSPtOMNcFr3jatQdGRtuNIfn/yR47nEGhoJ2DRVTc6mb2RjkV++qBzEnUNGhgY6Z
Wf7quaBMKJPO0pL5I13o7NVqNsF0KibEZ8pc8Todd/7/TmPO9S2WweGzZRmk0IJ6jEeaS80MjnLI
Ty2T78INdtSBfuBg+9jcNdzvh0196S4Cs5F/F8RbsPYjoL9ONiKL4/rbsa8wi9bQPr+CmGVgxwts
qQur17VHh7sqUPCjUGk4XRDa1E+vw6ikzOi62tKy1JmqFVWaxlm1WNqHxvmz+Ma07UabH5FEOWMy
70hWffepzmJFro7ZZ1aKndZPytjnsi4k4K0qIVJpAW9OOkT7le544MV7fBZDGoRTwvN4hIx+2ca9
1OTsF2pfULvVKOT2m295KBH4l/iUsmNzQKfpG/ADHZHrTDbKIxmuFJOKjxaKEOojRjChSYRd21rp
zxNiGhOHv5acLKnawb7QSgJLD8Q31DPTiG5LKKufiHMRTsBVuylgDrMmi8AmTYRlvqGSGJUZ0AkF
ltxOCQLYuHDoY5cyyUxSjYHZDdBJltUYamW+nxk7wMCNdiXQ+6tcZE/2TO3OyN6hqJrhfHIZUNzi
dGDUd58lB9sQaO2C4m5t7ggVQu1ORxM2pkDPL10W92qqEnu16N2Eu7tZBwCfls8M50D37Llzndk9
j/Jfdh0AqEjXFfVZTAPnlUBLKzAyqRlq5ykzDMA0FOh49kp1Vf6m3blhWYH4UtNOVw26RiG2/+/o
F8cx+/fH7Aa2oqMEJ9B+jqGdDw26aZweU/AQPj/1tDP6LNeayIbFg+rK94h8UJdaxSfH9bOJC42i
N6CJlq4P+0LlCMbmQKtjrwOwmm9Yw1vdEE8lkEhUKK2uddBncPvkJmrA9SgvE1NLG9f6nJ9XS5Z4
TrTGjpt+VYOn6oyniBs5Z4VJ2qSlZo6qwCAg8xEU+Prj5/SYuce01uVsfo1B3/LAA2LZOz8HdQVO
1BvZgk9kTHHHCse0qoAq4bgoRNO1ZiUnCd5m7vJ6R0AdfuaIc48SvpYssUBOqy8WtWxxS7LY4P1I
0c+x8ry5OlEmpXl1+BcFzXcuYyQqJgoGQNWBAN+YZ6FEJ5ZQjH7vObVBfwiPCsCOB0rvyfxecruG
QGCDp4VkKG33NlK4od//7DUpOj8RiZYPLKWwWYH75YwK70E3mIQRdeYYExtdUWR0izwOQH0G3qSZ
Ci8x7kINdUP/Vc0VuacJUwBZ0vk9yJigind5/9n/7WptkMgrTBPQgEZRfkmRgczVUO9hxr87ofyS
095FKQUgYJ8MWuw30YsfBjZfLFEowLhlm8VpZ8C0pDgaw2V+sSHR+LIwccgdlm/salQf1AnBsqpd
LkAP6mNUpx+5Fi7RDiJOEpo6Y7v1mJ3Jpkh48Ep6Zb/vdB9XKnj6wx2EZqMUZb31R7Qe2wpz2+r6
iNlQY7ja/6ogGwnbvuQ9gNRI0MBl+65veVX12bzVwl6YkRTOC5LdZOhufKYoi2bAVa/MAAoPkk3k
Vf/2gFxQi3BAc3mpxfEUBFxVh47CjniKKSUIn2yp6hNHQarO3oBkIFQAOpopqPmF2bvlDlcBkvhj
dc6iWZfBg6Heeb/d5GaSjgtR4RjT73eiJp3EEoA+wu3UYaShcMEdaWX27TYL89bcZjgQqZFR2R+8
75sfcmDmPcieFod9nBNkwslhERGGrcgoPLiqFCb0s5270an11liDWRe21bfOKCT3ON3p78GYxBuZ
krlHfLIRN8omfYpCkf71GCv0aKvyfPKkM2jJ0fhModR4rHvKqEcXRe7QIdT0EEHMU/K/Iq+mHnMO
78sQcgAXqJEU7PKErIMgko2HND7VraO8DgwBIB7d42i87rWGkHOZJXe9X1qNdVtR58W0gyOiuyqJ
upgMe0s/yCSCeViIhQ0leRcMGqY00GSiC8YlZgUuS49hoOab5U77SzcBGknTsmZSBJwDsgjnxNID
jfi5tpqBtImJO5D5hp1Yha6+7qXyC9Gn2jAgFDNCxFRMj2YlGI1txFApNEpk4ZTotloCr70k0aUp
y1dsmUusSx4KAWReTNT93DpnwYR8I+RvPGN5cZTcP7q/O9MQ8PA6aLhQOGSuCQ8raTCBdkjvNjeN
IJAqRF3AtYxtsYAecVhqMqgbrev62BENpHjxa8OGi3Q5V9bLlNgHxGz9oQcoHhREtt8DujtgEZFv
2rjp05wBTrkgbd6oZpmG47RTbjPeKCrCd3LUxmvtaYClq1a66dBFI8Ppu/mdZdyCC48o22Nvq5k2
3xRlswexkj++IewUlZcLVQPrspD/Nx3zf0nbpp8jg6GV+U4ZT24HYDzWC+0P+IxTPMba33Zt4ZOH
f2/13Bona3ASENLHCD8c6fyh+oQDWFlTmCRrXpliZ+A6DFksbgKcwdtF80jGRAsE5oz7wf6BbM16
Ho1hfHn6hOsgIPigMwiom8GYjJGW1xSCkzORC3anN2umwtqEIlQEQYzaBLH+nBMSK2iKqy/tTd34
5cyqEItQvIccwQnnSCUM0OtV5CTTjFJjMaQD1fvqbFZW4M8y4krZq9GBvUQHH7yfomtXMUZ/6t4a
dov02yr5Ecn7mAaY3cuiEVbMfHMLtUB7896WEXM6ujy7rpnOgcy5S86oPxC3P/mBioEdCnsdMN8C
xBE0SBI7+mueoDzjrWH3QHPDFy2TjhADF1Fx3+uLtoty9b6OPLGq6KN4/8nx+xRNdscEf5lmEag+
T79ZJIPa1JQiTJv2gGq07PB6Xk9sgx5yDXrtjtNkuri+aD4gJFhCBLQe4Yl/JpYf9owMHFYsGNkV
Rus7sq5ucxLAowFi6Ln9Bu7ENmxZ2Wi6YvYjl6+Ioqa5FvZBrx+9SpKT0KlLXmRQXult7NxIg3V+
CeKOGTRdoXSjTWgAFatH+VlD+a6GIYlcKlXCAmqjv/KPu90gf8gmlGd7IXqf43PJxnQ6EUBNAr2p
kXBkGnB+HGdMsaBC3d67MJjr2D95Zn5sjkjFzrS/QtPsuelSy7cdnRyoAXOmgLuSi8pHSGjVe1mC
iXQvBez8hylxBy9pptferuAvQFbGb4pqGLUuzCz9IzheeE3bQWLJpay6jrfA29pWGpR9YvDQeYU+
stIwXtv4hblAa7qFqAc02BIlgLSDBUr7SN/nsuCPjv3GKGZOY6Y9E47OBDUALD27Nlb7yegIYer3
saGCmkGpvp9S0nBXXjg1tg+GTvHj+Dv7I4Z0re/ca0KtfdNQAuYHLzg83P11A0Z/a+Q8WglPciaz
Y7ne2E+8kzm8zqpVLeGji7xRglxm/+VLQcrlgSjLwmdFVyklCVIunXNdUL4TDFqSG/kziQmHR9O6
xCmbb6NdLRMzsq19qWMYElnjVTHIH26xRrqWhudByja7XeSuGJxnvqkjAIGDvoDOCVoIg/+pr0xe
tKC1crpMgBlgptbUteO8y10forJWPqewU/Mmz/qXyKO1Syqydshhelt700Hu1y0ox9GJSADmcuhY
dWFYU+yryOQuYo3UY7rziuYxsQY1Sl3ouDU1cGIuV//J3JMoULMp5Tu4tvdxmjsBmq7Jb1NeNgEn
W9Gck7vFMar9sbZgX92LAmTDMfO2sILRremlkvVa8RbH6epbm+TolPH1BFK6fPE94h1ffR/VGl3j
h5IRyrby2g/RK6o9r/6tCTe0s9GpVlmo/4reMtnN1El7S77DNi7GJnklbiGNxzSPuCq89+AGzpHI
hOhwmHlIm7p2pZqAUQmlDiMQwiQazQAyKV7dNaTX7iTvl0vP7Dr2KpM/Z6vXz6Lm1YFfjGl7WrFy
C5QCVkMTcNc1kkWjrribaTv0xpZ3zBhMMYym17Of2DA2d0Yj685mU11/k/1Ka6wRBMv58w1DCa5t
H2Byj48zZyOeUca2+98flqrmb9SZIjgTHtjJ1MagP681HdH3ATOgS7ZuT5FJwjb1TZ4ePlCswnHI
hve+yf3E0+QJMNMAbOHuneC8jJjp2rxy0E1CbvY0+aPTAekGnuEUf78go/iV4UJD7O51mC6kFPFe
gpK61B8yo8BNQA4v2HvITjsrO6PsqqejC9LOSBg6Bt/WMMwtNCg1tjkKXRNGHfBXEdHbdxOn4orr
zP4Spm01iSx7eQzu6YVQQPCjJHb6ticwq8O/6Lz75OUhWbZdYe2EAmluFah5zmMkyFwSmP5OxLJv
NB3jcdXU7mI3zLoa0d9FX/tOAV1oaA9yWckQHMn+XVXdHtlgbQP/DyTfh9ecVpI2u3NbYER8TS+W
v0Llrd6YAzKnCGqzmtZaLhYHwxJ+FgvBd9/DIcdGE01kKzPjHpEMriH7QATNtWjsT6XFSgHqy8QY
NPOx4/IqRvhIwt4QJZzDTOyPbxdHmomYitnDJIXufKbs2EyXWHp6Y/fPIYhaE2MHS1AizzSqbSdf
JHcczUFti8GmB1k2yVrAXuT7bQYc9nS9ujcAKQKdlaw3fcCT4Kj87DZ2+VJk8euZeeKj024ruste
9CKxz0LHbCcDBpSIJkvUDry9kXHZ5kct+JRJuqEncoZCO1Ui2UV576Xkq2DGvPxRZKnDjOEDacP7
pmXKEp5C0q8mnyVz668wH23IQAm6kmUkAFhL9zX9ciDCfmhT5f+uwJPaO3X669ZqO2FzOupzkVZ+
K6caaL7BD7OCGmZvjA8YjtHGRjzLRZwwgQV1ANpHc3rbI/27tHJ/yrZIUUus7/dJ5eXx41lfaLHP
POi2IN437YD8nR3HlgOouY5hBiZyIxwDQo6Tplo/PYOETez8X25idsKai9zLmGMBLaw9heK6ZJR7
gFsnijzm0FfqOIwb44xATDkAWIRo6WlGW/4E9zcE5TZbgbDcyO1aFtWdb3cp9LNCvSHvQMKTnq9S
1u8JYnRK+a0Ms1Ez9TLOkWYPx24HiUspmQEOefxtO91uju000sVlhORkmhxP4LimZ+dy+X/8QuOQ
0My+L+lSR3tFTM64G2UpKZiLfOAVeJklSXKWmYRhM1fThKXOFQ8rLiWQQMqUELr9HiorNHcPqI+x
4E5/37+nBNMu2pZHBv0Y8MHcbrg22rKg5kwixDpZ5i9exLnrgoKDQaIOhUA4yQGDZYWMnFug0NWg
qtU1g2nBviEY93QbrP4KCgrtKvblwAqyenIS4G6kE/jzufb4s/84ifuYpVQ4FN1WdHbhwMi4VD0V
JGpor48g0lzO4A5R0tEg8AsHnpD1VTmpV4Yo+CUhGXaQX4ActMBmzVjyhxsYc5E4DZcr0+E0cX2E
ywRM/ZGbTf7wptPpzZNBPSerRXth/N3TvhTBkunxXEBPXTuUcrXfuhFCSLQDgakmNWCww7zqdGRa
TdSqokIWckzR6RO/ZhMAS1EBLbwHd3eJRLZNtsTTo/dCrsu4080uY8BQhaFCDjSkjJpr11YlTLgK
IxAquCFoQ4ttGHJ1loYiPCR85+wsha58+vN3Gd3jHhihXBLC86H4sV3Cbvb06k0knWtMxZ6GAwuz
gS/JnBQMfQggoPaEKMe9Iqit+C/Xnanp4z/5YFtgLh8KbqmD4vFlepTyso5+qOjduAKmd1IUThVv
OBFqQ/4x8EHPirWzzSlvIJG59ecBe/NDVd3RZCPYM5fS4QiIdxu+6DYleSCwZ9YbBR+8bZF8Lb74
JsTjwcxjn+4FzuG/ZdK8w9CSakCvgb/sS5J/QHQJZyE7MCmgS1wEyZvo9x7MPrNH6utul37NrCFb
HRlRxTHs2m8f7I4bL+A6VxILzkUjkHcv9tal+Hl91TAm/nA6tPWJoPVqn5U8jRceim/aQUj4sWX0
wnyLRwt02vUz60KYtqya++0UxaSAZ17Yg0d9IN7VOVDgmYHWQ/sqE/P/1rhaz/Whk0Ja0K9Uagzd
ShgJM5/ONYqs448kxEBUlB4oMnQ8/Zun3OAI9feXDEW2UOUKjSrOkrkBfC/YRH2VCraeKEhvqS0X
hTr6BSwwf1MmzCX5qVbuhjj7W7Q4qYzZad9BG4uEt89sc3gvwCX+1oZ4jITpPgnJjHW4NDTHghdR
9IpozziAxaLQxrOYB9Dh3iIe3GcUSZ3lcnP9J0xzRHsRs9uY3pIIDZrWLFNZgX0uRvsmdPDN2y7c
n6otRUC863NI/dFNXsGH6FiMiO298c7PHT6pcY10453r2AMH+m+RtN7GSFfEc1LS/0JXGgLBD1tC
BUunv3ihJALDNW8DIb3OBogcc6HU0piNo4ssFEnaamfL9D5R5nmjgI3pKzWs6mifdYJS1DiizUd2
dfjZI5gJmqkirisoTo9IgH0ZIVV2YyuzDII3UhWJjEKxzu9Uxi25VoAh5vdWKzLwvrpgAXRCpaGF
OvCL3qxSe6SPceD8GJQen9O4+qxYT43iBlZIKYVVxCIhFJzAzEGXb8jRBla48cDo83HGN+BP8fZy
7Mq5Voj9USQ69AsRFkAbmvOOgI1lBb0Q+NDmteO1vTbmRbvNtWMQMzXHVYwyV/qTjIJOtpVcosLu
2Wjz2P35MU3LRZqyFSKhW3EQk5GdwJT0kMuQEtlLbp91qkr3mLN+e0kf0doOQJ/m9e4zB6zGNNBF
ncHDyQBAcXqiTcmpbQm0sH3fa9ak7klT/NU3YquOLUmfFlC2ebLk4YpAkI3ii74CdpIeito6FN/4
V1jfMH67SRbgaAOmwE1Di8t1tlI7THV4YRF3Dq/axcnnAA0aNn3jksc1w52UB3UMoU7BykDjIkiv
CewHtxL74MolKHBdmYXmegwI/owLdKqxlufmL53WFxJpeAsi1xTh19n/rd4UrMqEEbTWl4P+76hF
3MbADZHPdBBWnmF4+mWMBHs3f+0WJ1qelXBxhcUY5nPkAg41P9I//4iHfxi6kF+hdZUoo3XQRYc+
PAVG8XxNWUdb9PibRN6dY9HCWfto4jhCuOniNExICaBP+WXtnauKChPCGC8dYo46VBUWEqsh1xaC
6rbBYP9ZW5F2D0m7Obu+2xDe8GZ7aCAvZbsK9zRw04w15xkJBdtY4aZuy3erGgJEtPQ6hz7hkrer
OLb1KGJhrGfH9f5DVufR1c76uPv9pBXc5lg7ZQMHaJNNqfgyNy0xMY7KpuSzDxXtWlw3RValq+bF
SvAx5plDNUaE42obXpvJvX3MBWnCyK9S7nMiuSoSWlTptloF7SS7RLeP3g9UJV75jhBfHtJoPkZt
XgiXKMHKI0r9cdTCAMBGwblCQy2++VFRGtujRniCO9FUZGj2r1jq5+hpLEXVqe08GUtqeu8dIO/2
d26p/pimNRWs7q+h5q8gMM0cUGxGTa7SANTMQMff9sHf6+J56BBduH4sXdrafaQfN1ij06M76bCF
p5UmuSU0xursa22QaU+83RfMqlj4Gj9OxFL4Ys49XUIDp/1FoZ34KALYN0l6ej/0Qe02sJFH9dHJ
vktb1YJ37hvk+LJiGnzNT8inuwvFIxAY5p8oIo8naIVfnACmQuwSXOvy+m7M8lofC0BNQOMkDK3b
00yqmLEfwZF6GyTvhNN0xHihaLW0OH4agB9fbHkP/QKg5ot7ZYA60y9Q8aGH2s8IqKDbE4embDS3
f0TuoUeGR7G7JoORqrXGbrz9i+YULu2E7ddZ5BB0v5FXuSLTuD2dJEhmQeWHcBDU8PIBJLBfUjOG
ZQtx9k+oqYwkWAZ8KYpw6Pt84rBzKBnUrzUtbJipocFPOEX66ULHRpp3hLEYLL/cO1282lcLL2Zt
OqQ0sJ+wMH1YnsVpFivbXoFsCdixM+51uhvCRfmM57gS30QB6n7Qx+j4hfNa319bBW4whQIUtNiQ
mlelLyT249ANKEvM89+XZ2CW5Xm2B1tzO7THszXnQUPFmEkJZ63evyw77Ghe1RJgKLTVQ5lAnEVa
/xZp3fnKGvTraArHtu1lKgx1kaGK4fgZ4frJ4HyNtJSZy35SRB3U/0YuEmNZIvLasEqqjtu0y0Ym
R4ZN8cJlTQQ3LW4DdkwxQ5hmh0ExumEQSzSHFvlwFwY73ur2mZGa/Hhe1Qy8nIkgCN68/5Rqv9Of
SMofCL0MoWH4onhVlmA+TIxzPdPmPxFK+Iul72OGhAVt/WU5JCSgX1LnWtw5abySNxI0wJkagzbo
72QwKeyRz5ZNqk2xhKZ/GXnLIC9OZlr+o18tIsvwah8wGVq/q1sMIrz0ymj3w7RUE4U2bOqdSXF7
I6Y8pdt2qdU1g+x1S8O7NAXBvOQczClN8bEbECdFGvYEnb7apDcHHso1YqxlW0kHFCWE/mQlKExJ
VYZzTtoFhqYctB0H+u09TtJQ8t80zHknc9BEPZM7Qslfmm+4LrhDr/By3lf/ewxddgSpSF+ujuou
bK2L0uN7nE+tJao6AYeTvN7vo609T6xFsWkVbDKg7hehFuDajbnX/oZvRzTHdqCPi9QVwvaYA8Re
zs9YNbd9/9QdR3GoMrzG/rTNNHQB7n5zxRvgZPwMyLQxJr3tUVglwt57xmOa0Cpka1QlK48aaw6M
3qgdKWYx45dzpOjV3jFsCllJLuiEXgoQrKI0+39SvaTbfwfGFQVZp3LpWhENqWW8kQsAYxgT6tiw
lhhDV9cPUyfeHlR3u+oSI/n/P0dvx0u09E6+I38Um5zjJEU6NEnxUZz8UeJ4W97G50xro2uiNpT9
k8kW8lQX5GsrukVmlIGhDlkF9ZQu1Yf3m1q+O3LJW7toCjPqPOv6gcl/693XsV5fBck54MyqZqJQ
NQ+LtVo+3dzYy80dhhdRdxu/0KEh3DsDLFJMmQLKw/IYv6r8jLG/7/UkTuHROIn4DoSaDaEqFGFI
Qc2uYQRwHqzeoV7+63WrWxmndLk2UcWQzooR8ywpgJgMOyJhPn/6Va4pZDwW1VYtv9PbCteZALRo
klXRNiC3bF0VC5nz9jOX7Mi+i4NnSmN3d30Wjek1SHTrX+wPPwlWbVHRyE3dfzclftnfu+owOEX4
4xwvHIKEODInW6I/Q5GIjGmbziBHXZefDt7YwClWr6zHRA486u61XDPA+LIrDxxc9k9THtG9yzr7
lbKBJ9LhN2beN2QKGs4Xr1hApuB/yyarz8Niu8Ap15RG9WRN66W4+d2PexUUGT6Qvij97mPGf4kX
IyLvP7H3vcM61BkFxvUIDrCTXT7Fl7McxdGJaKcfSpm3tLdA4qa75oW8W4bDboV9hXusCrJhcMbZ
ndNxpi55bYGaMIpOVlLBa+njYJlSR+N/X02OD96OQWG8UCqSKRh1l76bX9xILxYpTYhzGuPc7rk1
6McH2LSxJTuRVjJdDR0TBOg/t54Tm//cS6tL1qlK6YtNTR0m+MQcUjsFeof25t4PHcPcM5pz2bPf
HOi9qbh6x0ai8/1tXmmL8AZnyZ14K71IDUnZrhYIB6odm4kLgGGJA2cf5p8ZUe/5Kj4zX5kGLZLm
fuHhj1bL6Tf/KC+xkymK9Q/q2yizN09K3/C9At97PteZ1X6E/2agWwyEYzZMZl/nY+w7yjOCjqzh
waKM6Ho5ecxkNKQKd+VPRFn9zb+9z5TamHZjjJ4oPUyJACUqaFWpP5JrHfd711D7GCzQ0AEd6hJz
4MAUDm1GF6BICwT6Q1luF0LeU4AR45Dn6ra6LYAekPvquvn/go7F0Cs/x1lv3eMh4lv3Ztfq4Q5C
i+IP0ogshHqyaZB3W7/2LoWZybFb0uUNaLn6q2AXu44+HA3QbyQPpE13ZJpLLjm1+PuFSaHW9vBo
AKsmeOchhVHpUROuY9POXxbQlBTgSXc/DvjG1HzTyXRrpDvl63FqYh9PD6+8gZ0L79A24dXkqXli
uG2ixllnHxFu1VXbclxf6DI6FqsbsM7h5EOf5ZTuR89fLzeCXErxtA5kWkn9V9OIPryWaczK6heH
esuREjmQHW3gbeXgJuNdLKsNcybgJxNpmpLTRyjqeGjDv0k0/hvVHiWD8Atz9bICs0dijwtL6jAJ
fkijJsSbXXAEhfhaoa4AdurYlsbk28RUEFF/li/mbcYhJwv6i1vQ19jNfyzpSed73snBUZaagc/i
P40n5ZHEz7ZBUHXR9vHxw5kg86paXvH6NcRTwfZhIUneWQVBCfMfXqOlOFb013oVX4+ZoeQXXN/p
VSrnJbOZ2wTrTmM+WemXHR5n/VcmX8CGK/RDq6YdpPKnJB2M2ac9pwxCLD1InBv0SoCd4ImS3BAT
H+2fv125Pf1KCzQ9IR3DE7szAwlA0Y1op6AtgWIwEiiOq1Ld08mFWTL5XApL5GY+mpKt9Z/1GsZP
LSvvW4BZg44zo1E0CjcHnhyS1FUuVXj/kycxGw7RRJ1J+fr6BBOYP2p/u9Lh3ax+NzEqqtnt0l+i
1hiOiZyjvtB7ZtrK8xOt+0uiGhj/8c9HJUd2K/U4Gw4Xl7VwzZzgp/bXPO7nb/j+GHuUHROCHCRt
ilxmIsFxxxDZgFnC+hBluQaP7LpOVI/TU6/JcFZiui+8vcLCBHF2V6BzAzBC23+YVPV0ybjoNXkd
+QPwn3Vw+yoLOPzcmRyMet0rf/J4UlaFp4RrLNpTevS0UNZyGbGM+R2CGvA3KRknK48tSbqWryxZ
6XUmbXm8T2lfs1uWI797riklANjUGJCYFyRdAJsn+APeL4Gp+vg8xSHz8uQmp4kTYuMM9E+ooMRJ
r8iUa4B26WskOckDmKkBosT+USenmcncVVOsgviySpPd38daO2hY6iDYZr9hqIssmSbji0UymWku
SZ3CUUmxtTNR9i0HFsLyesF9vZodzxpVSVLNcflAnyDpzH7lNzqVOHVqG13y1AQrFERzH/5/1OPl
tRAvEXnjM2NxrGGogIFweCltCE/Fj2GdFTKzQRWvsvUaomBLH8f82Rh74W2awmfDpE3Q6wCNFI0Z
vHkH0oa/ZMlxXHVbWQww7RhiGZL5Rj/JnZT0/rglAduA2nyM7rCcsn0GoAclsfIO1/jDJB4uNZuw
Kq2w5/Sl9Xriz/5r90IEDT/oLD7+6dgt6docsOUl96lRCi+0BzllZOYck7WMb6JJWe5ig+eDd59n
h9o/x9MGRtZ5Myqc6z7eQX1J5tVB6dUax07BJx6zZP2wWuSI9yKtaqcAz9QaS7uTBXdM7qIL9E4a
QI8c+/o7HHu5oIwJgZnjR8tpBYcXErKxa/Cl0p/qNuFbYZkKP972eMoSRDUfzap+zQcvAF6dJOVP
soJvEyOEFZ3ZdN0DkE8WSSIUbcYAFvqJ51QVYvxvYCF4FupRMKu2y/U8RlKMcbGztXPLh/JVf6BK
8HZpQGBHt35kZ5H5snT7FcYICZ6yHbo8dVhxbswBfUv7l9B7FxjpMly7uzN+8tJ5OFNoV9Mjw8s+
sJsJdgNbKBUvEA+KdCYyB2kHEjfJt32WKrhcEEIXuLiddHgOkb+zFM7ayE6aVgXvFgs3vqbs6XYq
bx/KspeJ+XPfF6KG9WZn08ORApYAXHXzHFOwlc9BXVQg4342QnGjqj8JCjSp91BUEO3R7zC+Pmt5
yWiRjQX+Zc4TvY1YzKmH8D/KmI6vUHDCaH3mcIPUJTu5t3xRVeOX0E7BeDWWW6OWw49p2TuOs2c1
9xVxlu/8u2MDhaaIcEOxhuNxIJwBY3tgV+OJttYuA2eSFNwi9uiKHaeSMt+W8SqywRpVe5UPtDos
yZ9+xOvcQBA9QgC8tRpD77rEloOdjf/+MkEtb5rMldLfUuSPvb1G+dcQx14/6UkQnI6g1Fkt0RbE
ubQQ/SIle/K+7ZiVx5pCVFDKWchXoGATnrqlznIEk+BA33g9i6KrIjj1AOyJv5G/qAwleRRFJrDi
p3v9Utf6aQmQxnn3gtjLGpIjvwNJ6yPtn0eiIzGsVCsjcY8IHT32NhjS0hlflEBhXsZNGBC6XRrR
SMBjH0RBUxr98v9Joq1BwA+DBdkfMD+9GEMiiWunHLsmUr6ZG1W2QN3RUGHUr6V+zL0D+zoYvvkh
uL8MUcTlAnOjkxl0d/UrmxOFeQKNX3D9bU46oH4eDI+0AhatG3i1Q+ib9bZp/fLLDtXD6SfrPrw2
akDwapuGrWHtMiPpiBBh9p6xjI1GPlh79MdGPNmG+gS426sIabu0Y+/JoSw9VZGHZ3DwsTm2uHN6
wCiM/aTLSTm+Waf063HkTtAgeLGYJnC/MogF/NKerEPSoWvsnl7mS9VTc6FQJKq3GQXnSWl0vwoQ
gMVQZRKHbwCtvX2uW2B62NxccyfKX3KjclpfE3k00iuUXb3pmFDgCuq+xSEJlh/cxDgADoQL03Xp
N5NDlSWWj78mNhc7bQRmJoIyQVPI+jjU1dZJTCBZ+2/DZLk29Q6MbEXo/Tyo4pXyqzfeTIylmxQg
P+kMKSXaMMbToxU5wT4ygn9gj+zXlXPF2scuz51a6yC7YXwo/O5sW0+U854ON4twfkvffmR0vnfz
0Z1heGuYPwOTRyoa1DgBKN6s+owOLcJX8E8I88wpee1+xBIaWwJzpBHYOfj6cWavdTYHCpu0a6O6
9Muqto0P6nBylvbOSsnvn1gG9rD0YpwEE/r1eYi2pd3i7s9PMkuL+v4BRcvLMIWQXl6INQrQl0wY
v+8UPPLbD4Sy+EbCyokbBgzSHlSBIwShbZjeX4koHUKXHmEhztnlJd3yoiCxV86/Sao1x6RFnKZf
B/OsMMdIXtKlc8PLGq14Bi+a+feJsPyLThdO3wWmdh3e6Pqb2ByHwFSgEgDT0QbLVHXdBZ6ZaRXW
3JFJA6DAgMYerFcr2GL72UmvSwun50wt9mBrlNaoMpcFTXDfWdM4Beu//02PAWR7ptkLuCAQvTuA
QZMrtWaruMZfqkXQfSExHTVts7/gY3OEl2RPaW+VteYgPdyjEblPzApHm/tujZdc7rVL3ybAd+TY
n86VBXLTuDsL+7QqzyZNGySVtzoVzz0U3uwZ2o1Z3MfSxdJorSao117y1+yUJ/+V7875AflxjHY+
6I4fWKqJknKsYDDDQffS6WQcr2uCG9A1cgxAMTE8UdF976ad6T5iCGULqS5XDSBbMSSst6H0otAP
aOc5j1hNRPQOMyX0SXiiKTOfp9c2rNB6njoO1n1l8jP1edr5DK9zIgEGeg47z+wrzxPKcgzVGzEv
blfH2j1bSEH1SKPdTFd0c2CZR1luSTjJoggSz/ma2/L/Qfkv99JkxE9zHUrR6wooWIpVw4XWtcuN
igq24A5lIauig1oVz8zoSeBPxr89dHcl/GgdVLQ9GwRyvu0yS9cvFSUSsVm7TvgZ42pbukeWaaf+
2lXB0ULzFCncaoQujhDGuOrQBphvZgDrIh8zyBMWV3yV6v7Augz+BixJxS0i5CTK/1BtgvxBKpug
jCMcdHAyHtp4IVrRYS/YtuyBxL0rqSifkY+8F8SOpMs6QfwvQdZr62imKwW0Tv879IY0eiJ5sTwI
Fhx7rtd1y7PaQwKVIcfAxVfQsfo63FT+vhxMvSasfta8KUlJgwZkDwI9yfzsc3bz7ckRniwg0xII
YDMGxy16+3XD4tJ10u8LEizXvsLOwxKTFCLNp4sXPsURJjEEkh5ymuvsZU0f5weRzWCCX58vhf1e
XNZ63KUR2Cw69M+LWnzgHq8Z4KMFh2IStAoCq2YV7K1ajqECidEjhPtEMrMlGkboaR2D/ma8Fvmw
i88cHNqh9UGsgFg01A0aitK3dqsu+Rd/eop61+/q8b3c1KVBqlIfIss/m8VsOst2eDNmS5i9EeEq
2WWdVt5di0Z4W7LQp7u8rrCTBGKM+TSRDmYytlB2Z8ueImRnSns/i693QB4YFZwVZEzK7GintN2S
XMM7MCucY5ttbInAZhQvOw42XyFjVPjeyC7MFgyYsr5OhUikz3go6+yKQF+kATyOe4txWMfs7NNl
T/gLbgiHRkXIWjNlmWB5ODXUNdzSKidBpmjwEW2NSCpePk2RzqtjGgrfqiXOn7P/RgxJRzPiZVoK
Ctq0lj1ZJ/T+bn+0OthEZhdlaFilKXot2Gi5o4N5iT+EIK4ufVFwWUBeL4z/nJ5RjAe+rlTN+bQD
oimg415PP2e7v516jW0Ylj8HLEtohgTdmYQXMJwyYZjLH7pwABIlohA+rMhyMA4oXmOaX1zTTk4g
Jrws2WWqDj3VHnfgYjEDWqTPY58ygFebG6p87c+U0GGAOsyxyfWpMq1zXMurxAR5obvyxvLzcgRM
esvCxKxU8vi3M+MmENjVSScBu5y4qcHv2OMnjSuXIoQYw5mMlKYI6OE9DMB5Kec/zknOzNNSdEX3
geNxrCsKvsXLnnkjKIBCjBieThjf2DOAGkt7MCb3SW49fF3cEanR4ZTiPQ0Cu9GpgjVGoNt6Uueh
IEivJMLu+2edeOk+T6uY4y4gxzp0PuPDGkXFDV17VNq8DJvCN0r54xJaDVa+q4dqi9p9KPE+HnlE
3ngKg0gCi5xVHckKmo+ihKxqw9+/3Wjg6pKDa895r5n6bg8+rt8mL4Uv70PIw5/Sp/LN0PxYqax8
7rv0rLzEUUC9544bpr6xSXazE3+lpRyEE1eSIsCxDCBeFkPuzd8YtITM+7XOTNl2LMHQLgimZHnW
nkb9oAxEa3tAFdyIGE0Lt5DQk0QmGrPCY9FN6lUU0HkXdD6E296JFpZF82wC5lvXCIdeoYTtK4IA
DsINKEZkCeUG4JQeBQhktH9hjAxnwEqhsY0JCdipWkx5c5HvcxtmEkjT17Cxsr4yI+0R4BaQ+M1F
Fs9/IVnnVQuT3Qf9sMgFQmCoIcWsA9ppHACXkTmrEniEh7JxgRdzX7AS4fRzAYkqDvu7MIQ7560D
LEfebR+TyZDIVbKGjzH6XJg+8vz3r9tMKE4y0h/cnCYpJIJSgOt6hI8DN9Z6nDBjVLOuncVd8T90
q9rYa+Ild7JCoqKnet7I2vemRGHT12sGTLWuYCVVazIZzqpjVuqpCQ22MCyCfomIn8X0qFLR5hqy
AQuIBejUnOFlstzHsjGLY/HCeueZcPbdxSdY/hZCeHBmKpsJw1yJxI88ritWg0AsgtcJKRZXhRTh
/M/UPkn/7t9Bvyb0wpQV1IxIG0bKaAytufcAJAB5K+R5APYwtvIZaKYMtzxOU+fWlrTW/04Ev5tQ
NYfW9gdgrNOTTvjPhLcdwRuhNrnzlUulIQCQ4AURMSbXmAo1x1jYBGYVrtxIr4LNqA7PnsgeLVwJ
/Y26GD4eWT4YKqvfP+RGqmF0P4GKI6hUgFonmuF7rsltKJqC3pjxhS/V0SM7cAMPbt+ikWxSHi99
9UfEa2AfCAbKR59xVYVah5Up5aDQxINR3TMxkR02k1rW0f7qrg6bO9qj8J1hZrNe122bD0btvqpP
135oyo5pCxyQH8gKNVlxtjlKz9ca3q7nXr6JaMgtC0JjKdI6OmbF2pfzg3pYl3CVmtgmA/eiSpfW
0bvhCifcu369qLHLaP4fgel+3y/DjSKBGeSXwTKY+aIzYcQEgHUGPi1p3y25FVHYymOwrxstLTf3
oMHMMxWo7/TqlJ4l4oBAQuS60ztz5qjt44eeZ7HRJ75F9Zju2jkN7gjQKzseQbIJfBMoP1SzV+us
MITYsYvQON7ZR2FbpyVbd5OAq+yDWFsfoGPKPQQMxRdglLQCAVXkkuTIyob695WhjkR5hRreLJu+
AjfuE6onYzJ1zmL0B8fmahNxUrjWMpC83pD2+0Bzn62axMMUGtmuuOJ3IrWCWEL0+HdGu1kMds+a
LEc/4vNTLs7Tm3pxP6YyO0PRP+Q2GLxU3Y3MRcBGvPy7FBdIMRs9Ibgm7WQUJAO/YPAoKdkqZsvk
sY0sPS+RZR2e4h0WuQiw1kRJLoxt2TUc+XhFWDwpyUKe3VPXF7ZPPIRTtmPwYfiiEm2hOX5ErxFg
BGlKzBWmtT7OHReMom1U0928KYVFeNqtCskunW57XUPuDQylFrfb+BP1fwcjGidqRdYEKYCafJ0v
pHNI3I1YEHjk9HmncrHsNBav1XZfDxS1iuxMdaCfl9pSOZHADRuGS+ZlQY0ksKOu38GsY+ZEEBK0
C4bvjQtIhXkvWKtv4dgRfLfekYySIOgcfVTzQvB7fW47ZqPgf1kpeo3HdWX7oS60n59UzIQgJqYo
499/hqqut9Efr3SKNp9n44VSYTjAQzzeChxYM+2tp49r6Kz+CEdgY7YL+fMTdzqUt3ZuXwC7S4W5
ZiwLvJgtEhLpPYkTqXgEzD+LM8U8G0PUHcvsEIRNJQQtd0X6P9mnXbjShMEvf4r9wnqPPVhUWKhI
BnilB5XTtHK7EBYlk/sMYCftyL8RGd4kbvqF8Iz3w2Z1hubh00g246nGravkDT8V+DXswbzHbcXg
DWoxkO7/tbXm4ZnysCRSjHT9DNSCZ4heQ0Wmil12JmXxmOEKcsqzGdMYzwUmmECZ6nm9b7SxmRnl
eZU0JtTrQkKIQgL+9WbEVJBAoNqrikAvUI2uqbPpmXOatpQUdgrnMa73eB4PE2NKSjUBqnTGgt1g
1QbFcVvnmAKguoWuvxC2x9WWec6LXzxn4GTBQVc6EqrK5TTDoC9JvMWjFtkfkeeE1ucwglxZpyfw
pvjZ16BQf/N51X3M47gE9O4y9Q18k7uKFfVKPYT27Buk2t/bjNy2N4yunDy6qNWteSQpaNls132G
0wXn3mQwAc72y4M3ftgUYTfJ+15FUuPycZR0q3wJVmHoUObI4Ny1BB0ZzSRAHcWatZ7ZwS8IjPgr
rJyfUF2kM4jb4b2P7dpvfHLmQrFfoeiVwj++5/8qyh64Px28sj+dqupzMsbz3dvsMdV6zTuxQSVv
1oSEYOapkEIZ4SHHTOJfhM4szH+dSIZoNm1YDQ1vYAp1EZQKlrqANGdGOExvWwbhO/YyNGv8xIYZ
tVLujJLnw6deUXk1Tqw8/SmXXTBMuQfy4IHPoY+bQe/nRRGlKF0/9KGa4ZJyPD5kVU9jXWyCI1O7
QoPKhEpje4dkftRk722ElIqKz9ibrQrvkenS0RNNGKclSrdX625qtUGf45ql3MWMu9dSOL40q9WU
EQmLopjrVIfebYAjqWgwAicjpye42znUXt2kcVu269pUCTYgCrIoobhqYMi7pCtDQud6rV2nhLQp
MfEsQnFlof8m+7AEWrhuUXQTMh+FzSx6VLBzKtbu8IhbROAyWC55WzYAEaV8lK9HgvVMVq3kH23S
BNd40+d6/tbb+k/UHzzTafOAQbkDDhLK5zqhDKro7ZCrYKEpGG/irwWF4p9dezuulwPtyfBQPFd9
Xtn2mz1gAOk9m04mqXPXCkmz8n63RxMoc9y3CDBHgHIdcCGL68uRJbT27rJh5vvRhvZUSAXjTk2p
f2bmcggo4y+UvULm4zKeh+axy/NE++TytIDUEsMIh4FwWApctuzX33q0Jv2WL+AGl7DTVCl18JIs
r6dqlOYG6jHy2GHeWGUDRI+3pJI/4mpCujD1we2LT8/SW/guNcOTimxWjni+nAdjEEblYd/yOSMC
UB9tg6El1uh/dZmk/YbpARGn+1pKvSE8J0/XjZfSOb0X9nk1YCzxWgwp0c+TaYIhK6+WegkX7DCw
JSYCtlIhYlneujtsra90ilg/MrJfTzTA9autNWFaFPqXeeXjwbeR3Xf4YWFSu9lSsYPQGa+HpSzd
YNmOPFYlu/ufqSic73J3LW7OlS2ECARXDzsyFjlNl/DdIVawZUZUeP62xv+RaxBy9IoRokAXYt5v
qFMqFspzScOWO9HA1I6jkG7iYLcCVS+JgQf3KFgxnsNwczcPDehqaMIUt/iotA2sqqnTTJ1Syxqj
ALT+UmjFJxywYiqKth02zD3A/Vxf/p46tdoQ0/kuDYZzEwvxi6sc7D0okDPHI4Vg4E/Gka2DqXnn
MhJJsZCisQatkdYhND+ZO8cQXrw3FC5cMwsZCpyVfbmHRaHRBOhLNy6fP2S01x8vLBJRqf7D0beu
LIOtf3mVQNyNtYYydrkDdfUAjcee7P6UGjix4AaKDHvjEmnkM1t3ZvGffZHDb8WgWkFsRO71X8f7
E1Y026ADektmFHmxi0QcCQ+JOho9gnaWLUp4FkBOnJbFnd606iF7syxmNJ3IwgJtQAJyN7J/kLQ2
9v05s7phaoH69g0+W9PRBK1Sg8U30aGmn+8TFdsqHw197wvfxhtEt8nquHBSNb705ZFPwtvFNHbN
kYnS013cxf9tfrKzpvGqXYM4N3tc6QMw916KoA7fDBLz6eBkd90Lf4vKmFVdtq7eUgbqg9ciYo0G
DvRaUZl9f1IijPJ/O+YaK7RkJpXUDRmaBMOvyP8WSyaAoeAgEV+zuuAtn81Utj2m1eqD/TvaT587
Da7Y6IrMhI9ZsvKexOllYR7I+U6E29gTKp+0LP/iNtXhZIdYs6U1H3fmqliUmDB/HACLGa1eTQEW
fkzM38MBaCWxRpDfU3/uWCN7LEWPK/pNqjl1qIsZwO9OTAuQghvkXvdRnMm8RP+UfdUWOERSl02V
9eVg5b3xzcEf/maHPI3WNMoex2WwSo4cJ168rNKY1wjzHz1syDP2Gh4a3V9bXGvWZa05v22mocYQ
viCNAbPudNdpJ718VW0yqQ9UCkYrxOFfut1cLoA8rzdPc37DWsl8NRVBhcWd48IXiPVikzsX2RDC
8rTDXFZowlhthYaAiRzkEdrOe0X7XQY+XTVG5p0+AkmBVqcTUvC1sVQJu0otphmZVCgUkjAEm8yJ
6qxlFqaEd9/Gfq/Vgs4cHSkxzWcf5nE2ruWTt+Dcgh6kPOOjk4MBfklO4LuI31DE+Nw62wEbH6T7
kL9bVnjTLhVrymwjw8dbXgvi3DpMgMQD2GQM6oqj507x6uVPsNi1n+k9iX1cCxIty0zW36toVh/a
uPKVITjz+npmDV5WA0xulF3Vx3leJ8rmYkH/riRysnf8YU4q0X7yd6Hw39LyVCIMpo0/ndpBbCvc
wpuzQYWd57Oud8gXmtv3Ws8FHesC+qjNkAT5pJhNg+Z880Y7OgnJ09dNRhUJVOxr+HS+OmZ/7X35
Er1MqcYMXCqtH4lw7vhkQZGGU6QQDQ6hqwkd2RABNs9GnRlCIowbcjNARUJPvWy/oAi9abridYj8
CE0NfodQVm9sWfmM3qGyZeYDVle+vzy+ltUtzHkoTul4DOm/7zQJBg434ZrSIGBe3yMXe91fFks9
Z/HdgsPzQ5eJrgCMnWK7sy/pAKEKSSjZjLk+S7lQ/4CaIvZHKTtZxxMCWANtBXWDSqzB4Bt1OS+1
0nrTRSLyRPUbRONk8SHgQssIcLhiW4tr0fF8Vn8JxRqjpfniwGjkFiAzFuBNjDGX0necRhFXzbok
E7p8WXt1jQsMW8vyKhXVYqpyiv5O6uKrd4iP8in7djVbr3hL5O7w6JmAMO9u24UMmXHCSXhdeJvI
NgRyBS0G8EcVzVNDn7AXiNhVQYEA7HoNukepvp0V7NGU3W9rj0mPGPmUYb/JKAFuo4rj76yqqHIg
SqKkdpEwfCi4BmfdKGxtLRH5Xdk54x9ab957HzZqQqliwnsVYfSmP4Naea/VzCnqojzwjNtPUTpm
6/vrQvWqTbO+oF4NkJ23xjQ+3zVG87Y9UT6+BboBvpmq8WeeZr/FlvbfGWZurPKMUlXUJ5DeT3+w
EznIQivvy6mspIgLuLAZFQ2D7vE9CN3kif6+r1TmLN7pZnVmP/W1Opgtlea6+GEIIZuJd2dVs4m7
ezSWeXgGpG1lLZ3b7Fzm1JpzwfZpZCFq7CmjCxQ6Wwy8BSeKLVOpjB3vOybr0+EQIKNULaloypMk
jUurWmQFxrGPpM/qwHRXgNh1vQHt0JCUp8Ew4hGJlCL1651VRK75j2V6FD/4YyMnPLQ3w50trDxX
oPZqzMaZLI05v/1qQHWDbIFMzk4IGJJ1yTR+2DOiGcWwLdyR4RoIitSmnOJXIMw6Xoujru/73uX/
SyjC0yfrEKm2VBxx4XDcV/le3SHMOygUMljFKC/g7w1W1yXkNY9A+OxDwbS1jboHRDrwzGzC6Fkf
34cS7SSLq9Sna7eoz9CTGrVoi3GPfYzZApkPtEBT6DOh6uP2rW1bAxMYbzNSJ4emFlNKTj0oBi/J
hsYnvY5wJC26V7OaEW3ISris9HTtE7NWlmEgKXBakU3uBjMxknyC5Tf3lLJxlxFpeCoQ6vIKtpX3
5tYevnCuWrYAv8XQRBvWfXBNea7CD2e+m9BkTDixpqZdu9Tmny9PzLR0m2TemSIUE8lZMVHFTgpu
aEn1AZ7iej5774tZezML+vtX1rsWmdoGHR5xNbYUBxBpTHpRsdPGuow+RKJYra4caU/BkOX2MArS
9oyxXqmnxcYOi5I2oaVFf8ziHwnSfeQpir3IdzHIE2KBd3Y9DznTPGCNx5+/71P69K1ZxuZImcSv
uhUnDY5FnyN4MKYuXU7WzYh5Fd1Qlx+Jdsm7kZ9chWkJZk1RNvkDGqEP5RDpUg3uIwuo1NDKy5go
EDFZ5rd3nuOTqYyHuR//9RE9iQyp5XhlRx+0YF4ucqEs7opzP3t6P5H/admeOnTl1ni6ZdcE7/ef
+tabg8GqmBJC464rxF4SF2VvKqafhcvAt490ZW8aKFafVOpZjlyLE0qcgyMeyfUcTTBmslNSsV0t
hbGijAxsNMj14X7snQT4iteoGSeOO6t1+04QzRHbyhBJa3lNb3ANzpbIsegwjyxytw0wPQp78TES
/+/oRBJzPj2YJEfSWRO2f72584tnH9WZVmo91Uh8BM5NJejer5CWdroTcJE+5Z4URzVh1GA4lvX/
g3IL+2zIgPQW03CnXx9HaeeNfMlZgBGQW/YcQ93+vqpSLF4m+p7NhMA1bj1VG1eSIomJK8BTwa2x
f/KBm/PiSYiOC7cQ3kNjOC3m9pGl7WTtKzwKqN+NbgsCy889IxmUZS2oKd+fcq8l5iEBA88o/Vwt
8jCj+vqTmhj15LMtPf3RweNxct1sS0dO8fL5a4odb4kWFBUvQQBMxQn1WiXJv9H0O5JT+o2TrwlP
vrNIrhphjHp0PJ/2IDWKtK4Boqj0Vc5Fra11TYoPJ04sCkBLsV0vQCmR+n+aC83GNhrERIFQyNuS
Pyc00mOpeYA+MBvPe1AIFMEmZgfsI/hNm4CnrsICAgI4lrXZL9Jfe1H3P0JjidpGSTvi26V9uJyd
KkWXd4yYdwOB1goEZchORWD5R0WBIBmrdp1nNvg/kgbu+j2X7MPXSaS8LyNgBLCWC+gOGMEm3iM7
tZEqXFO7WU3cytrAMebHIepv4fmaTw/0NzRoHkO7r0OEXB+ceIV3Y8XFPo+V1yFtvBowFJzIjQi9
w8sHwn09t8FgyVXwX4nJitBtJBYKcNNCbGETju5DyZRqlkFcBBoVw4T9ALg347YNeOe/cIVBJ927
uQYadbctNV+aTXaaWsjR9+9NNJZzjeR6qx81RCNDeQhWbrHfGxWZ6k920QLUdKH0Xzul+K7VkDFM
nMPZ+X8PMyGm/c1dNrP1blrRwDFb9OSV0wrmfen0FUraIWBLEoQeMDVeeujKMiSiMcFdMeKHHRbx
/d8EoQ1hqrQn+nk85Js4LgkpHO1dJCqM9O7l049zxH4CjnmBedVFXrY196ppWO17yZ+wYvOX3aVx
pKrDm5/YYGKCWswTeIQDBa4jNyZpW4TSMBR/PqH9sU2xqm40lZ+KLVcPUzBav8nwzgFZ45DyclVC
flXmETcu1FPxi+X/k8oXpyyU4botaH/qfwG3nxSXKUNNAm+wi1bX3CII3547XsLgyGyvB9LOThXN
T2zKNinfrKOSfU9iQ60EUcibk9QMvWrneVih+/WmSXWWu2trLWl4szx6/VLdmFChcP4364p+DxdO
XPNR2tApr5qx5FmLe3fnuSFgifhhHL3/zG9ymv2vXqt9VRbMJQ3usWcUZ0FKb25pFAkx5dJyjfYz
fxVNLDHbrc+tcTczdY2+QVdu+dtwsd8fVVCZuyqmwXxkOwozSBqo7OiG2JJzMwlTrUuw9T1bF7vJ
YsF5MGPDCPxmw1i2vd5J0NYlV6SepGoUrJh+x6isuWmpfG4QQ3DBxHlRJFAnzopcEmgvBVc9joOJ
C7MVHD7NA20/+7ZSrN4CpQd2be8hEUhi1xZz92MXRi1khN5T0Ig2SmtN7G1sKxF3UWuhj5KG+yc5
+Kmh0sBkW91lr2bJ4YzEfD4w7RM9IJrwant4ji0NIZRtD41MWHJugcdtpMisBQv5oI+MB8xryAr6
qr8+1ZEi72aUApcsnOnWpskkuGv2PgUPa1usv3k569B1aFMb2L6mELXkOWOnqyNAGlR0AJgqudF5
abzKnj7AyDtGW0ivoZTtj0oSbPyTNgYeI5+orUNRH8+60izsmpNbtVs/1hNWYNjPRp3qq20d5FCD
lBLs/Z/melZ3oCRgb0vtXHdEaYdHqnyqszKtkE12a/rhOgXnSwixNUa8ciEn67XjMVJYapm7WBzC
yEcgvOTYkYkPsLTlG1ojHKq8wBHLw08BvHNjyM0+c+PVY3pCadzfQwCN0HuszvZ3b3wtOGMTKJz/
NpnFy6s97MspeVDVurP1oOBoxhax0aruIzATL0azOd14GxdUGlULCfDWfNWLCDLhFH9ma1TxSx4G
kL3wSsEr1EiXnXDh4QGyBwyhd1g7LDF0SiDV8MLPuXnahZcFdJPK76PK2JBku4qDEiI3MwG9MHDA
RViJT3qW/QEZNfnffXEt4bHyYGw0d8TFd4GAyg3fejO53eDGQQ8mCUukgwiCjWrFgTG8/PX93red
Wvwk4ZmrOuSyZ1XXinutaR4Bf3mO9KcEmvfOlsy4ZYAVSQJSirsItlC9AqdAnZMezJbrIYgKsViV
VEO/sPJOkTM5XqS8X3VXk0r0WlIq6+GWhrXHaDI8UtOFMpPTVFpxO/1SviyfWEQnpYiUrzgwLhOi
K6AnCu32ovbdO12k/ygkx3G/4Ya/FJ47p/K5pyEVWckNhZBwiSaiwq9PPaHJuY262dN9gnyaBh5U
KHszbdH2pEk09cwjwTMwDjcMm0A7Ti+Oo7F4+/rqVV0Bvd3/9aVewReQESynaF93dyNPNzwMpt80
MAyWlg0NXRATv7FNSzgiu1ykjH1bXRtqUEXTTU42Qu5bhw2C5guYY9zlJrFJuTfuOST8drhXLkRX
GrvqHWWHODq9iZ1YDEIaNjK+rt6xawrF7/uHHn9BJTlSJXIZVSJboQOzeN5e327ci5GJSy0SM6sS
dP4wFyqswu0PsCaH5gfjdqKf38nxLBdVnhrc1oVmkweZIR5oOaRid1R2mgFBQbZ/UnNWpKAxY4Gq
blaQn1vnnU+5ZFvIaT/Ey2HerxsD/YQ6VEl69qubLVO9kLFdXBlzLhq/GxztFTurQrZe8bQ6w252
cF78LvaLDJjyxxFLhBZOX3j2BxYXFP30oBFl8TTcDWI0zcSMGTv7WPwHI63+MG6h7MKeMvJES4iB
pRyzLH990Q5Bg7hL/4T+GLfGSG69FJKnzgwfiJrZnnkhI5TAdhLcCa8NtkLJvRzToBPHBbnlPEMb
ngHerHEuDgFyh5NPHz4HYuqiRXM1uabFIYtur0rNNkrL0d1KouD+CAXyCC3akvfEtem/ycE9mdl1
GSXDrDVXz25BhQlwH0JK1FZgs8Nf1Bs4o4Oj8WI99RWfEQkseECfzRc9DhLvp3YhlYmvN2H7DhOH
Zn8sNdvq9J8buXToZyz+0P1GaqUutRnf5GNo2zFRSn+04ZDLd+IiDLSzXDjQdlhm1wO681KC9mZT
nfF5VvAMWvLxe4Ood4W7DLrGnNWAa4bR0raTLxHyApVChDp9VNE9Kk5g641QqaTRyoUg5fXw/fPY
iC3eEDJTu9JR3bNcb2JkkrSwfOBNNGXPo3pnL7sBNqAJ8RfF7HpnBwtm1FrNNLwepftTsxvk1iKJ
Tn6cQfgWaiyB3jTTnLfDKgn+h8UVC1ygjuVGLjZv/iAnqlugoiNFnlxRhRnWNAMvtabMMkENbwwn
vBB2zvlhGzLX+r462xol4IAsyTaxawQ6OAgwF/orWIoKeL8G+TSiozpgWep9qxLPEjF2qeJMFh93
Nl6vH4+CYWIkH6FvMMw9YxKe0vwg0iFTeJUaWSmoMDYRoClCi5Ch3ykzg0sMgsn/tWj4aAu9b2L6
cL+kphz9r5l57Eto700BfPuUAhVYMbEUd8qsAIdlOxt+XO49hMAJFzePPQ8YofmV/+S47YY3plw4
yWyfmnEAT/bGxfZWSsIjY5SEr52q+L7Ic5dUoRUMU9B/h07g6Xnzksd7CcSX5palPDcwN+7VafIi
+WeaCngiSNbEDJCKXVnExGy9beKqL9jCb+MvhdtQQaT/n4VldxkctPAu5FOGE6b7xUS4nU832hvx
/qq9BWYxgWUDg/ZQOM1YJngojObJtL08P2B7QczY4uremcNgI1aAlXVW1+dHMWoWs/k9DnNLXV52
r9NiTCYpP3uoMNRZizvnoT5Ff0NPKfLMXPDSh553IoIyf/nA1te2cvlCWo8MfS8APXUyjOYpDw+J
rnqE7Embxo8pq9+ORk6dv1Nub83xQg5q1h+CFTmnytuBkF4tIqHP9BGuGF4KHrpkmH4XYr2tbB6f
A8kFE25j6scDd2mnEJGWznu2yjfqSSkapCN7L7WHHjnynVLAfgINgJg/Xq75rqTPrO5WesN6BFBE
Mq5SXCwkamVRUke70oJb3UlgFY/6/A2P75NJYxxPwQy6Mx9RgZq0HVXQhuepNamWHdTZccYdgjpv
L3P3vHFqOjaxPZMyOZo7+edSOmulhtKcMLcblKvFoj9ilGgVgs5n8N88KWMPxc+uyKntt6LPqHQq
CNj+ZiyDWBdy3hplTiwV2JCDJDBp43wQ00o7nRtWz8VPm/jhif3aMZJBXNn3Qzx0+j3fuTNmRQaM
LterI41OOnACJaI1CtzZN7S/T3l4YpLowuSOc2XXgI0oRoZbOBncpD0E9qWyZfpiq+8AHhGbp7X5
Or5c5n/PrY2JEKhDW4dvYP583Yx37quMlndY0cBU6gmFl9vBcyiHo/AGOKpJOKNRjA+XjAdSeoCV
XWEMIHeibE3SJw/z+f+bYln55MK+vnTV4WPLaKwl0MDKs6NUjqmWVp2Nu6i/8Lr2lD/7IJbTZGQR
g1EcnuD4og7hIfsbjl5WSWFrQBX1GdV0U/xfQC5yTnJ9LLsrahCxR8MtXAETg7iXPxiFdmEzILdf
AASkY3auec9G1zmgay5OFH6sabZAEDwPIn0qe+osnn7zY3L2L0uM0ZE64yZobapcM5x4d4cOyxTV
dx9mIpBrrjP5jHbLW37ot2bz/+AaEHdizJf5Ct4XwTyOleMd7wNdLYxecXxDWDztSnyBBcguFVhP
WMNKBqLF8w5QwLLra1GmWuPEDS/0PNZWKcoY7oPO8ZdBS4up1GEHC4xBe6JhPVpdiynuunFwb3oZ
V+fWugyDMrIqxs2kvjnf9E10tuW1Q5wPbVoYfj6gsUWBsaOdM5uyzc8Ndh/CZuIwbvc8LHZFIGFd
1O59xq+MRO6HtmjcIgkPLVbIDcr+WMjtE3T3QzRsd9Il7M0CeYt+2D7stWzKPSn34183ZcZGIntA
lI7P2QqWLPPHa90dZDMg0/tmtk62CUvoPosycZTNhtgb+vnaEI3EcUg1pQGILLGv2WFAG8iwt57R
rP6pvv+7MWVr03Xcdum7uHcPMjTSlF+9X34lk/1gxzDv4Cg5KivJIGZVSMPbwRFrIRR9eCmBUUXy
oYoQMFgD4MlxU1ykjOfYJsdFTgfYUpQTcNrWTIL9giphXeYbi/vPc+ezpQ4pqXUYzu0ADAz604pG
iZjnlQa4qJUDddaF3RJSOPS/0cbyP6sLYTUN75jkEguHkQf33i/y2vNqyLXKJbtte69Vf3JMOdBW
uCMLodlE0VMpo7/x1blEmpHpooyRH1XQMR/WI+z5H4alzklae0iZxePc0vEJmySKPBF28xWRwvg2
U7uyJoLFmBUZXol+bCBHJDXNcuH7C8oEr64jkgmNq63vFhveDKodJ66A1NUZVa7E6PL42i/i9H05
m1BvnMKCECc2KIh9JJyd2VcPiY5qEZKxjhDoh8z+4vn2pzzo5NTuMNjc3R8gwEF2EWvuK+KWYetT
xqM4/j17sUYXdnFv7WOLmZzz8566VFjQqcSjzRPQ6JiW4RGNJwWyLcC8/tyKUbMdu7+kuj68eKDg
rtkHryZmmtwjWAavFvobpgRvNpVsMpVu/6Ls6vSw3iCZw6CHRpLqVGQ+HpcceSETQIHSuYPhmrt1
bNM0DyKTlst7LmYlurO9Kwwdq+1AYOsEmhI3aQ0/1nZryqR8CGanL4g8p1KDtC3G1s15XvluRbMU
BzsCQNUHp7eF3wPGx0x7kyrPzsicJlDS2HzY107VRV1noGeJ3DkHI1ohwYev94CF7FKK8v/Av8nJ
sGSkGCuHtr3+6xE9VkUF5IbS65OWWJCbkjeZgPWUXkr/1ZfTkVM3JAhE3cjAfcI1goHe5RjJMUw5
wDv5JXjHiwgRWiX/oEkClCLy8lrmtMEKlJ9VBMXAU1P3TbLn7h8IDmai9cjo8Pv2OPTFE7HoRF99
t5fJ/dR+Bb6ESIG4Ph/02ORmCON7e5nOs97uigqbF/YjXPkxa0RpZSa3hCYm8bOBl9kutnREOSxu
99Rxi+WdhzmxY7vfqGNMw9NmGLTLLKibr/0KFL65Own0mdYhH5hNfM7NrrFpFCrxeNGF4zRVQ3UH
ktUfLWr4YfGfiJApxMqxinSykfMw6KghBpqNgZx5YBIuFdxYE+jMCVpupOirVWsJBeiR7Na1NkR8
YWXIDTsx2JRFrdiHXktr6KwW9OedFYxt2FUwnAR2tBItICRD9ZwIl1UHpWeCfeSLjGYf6NuDGIZK
JNlQL0vAvLSqTlgJCVlnx6qy3+jtjqixWHcjg1cjJV5ra85MC2+B181QyYoPWAbw6CGHLeRYRY90
IThLcn0HFGXo5jTRwSk6RW5Dadjrmz8T57AqMzNR0KU2v82dri6D0cv58gexpyE0ugwfdrwRhJTL
X+Q/KYSPP4dmJwRdUNiMBjxnWvKAeXwycDzV0pw6a0tKEycQy4ywDRReRLVt7/wD4MMDrrXqnsFS
m9X3xwrx653Z8VUi4FK4yPwJtMHjaEdqbah24lvojoxdMSVyCuEPMAJh1/F5gOLMTiFM1drpu7fu
oybN41m0ASXsf9uKEeKVMofbbY7MN2iRMaZoqtpls4R2CGWpto8ZdygAayRZyy128KpHjGPVqKni
e8Gv9uGDYkyH1Eji8MJvy9bLKqK8LgQO5qrXDztR1jAqBhwNS1VMi/Bgo+q+HCUOPFo0/jw4bf7J
ocdIkgxzY1YiPnr6wKzsxqywBbYgVRIS3ccPTjZf6zP9/N6f+oTlTGgim9FkQGD5XMI1eD7JLEB+
TAfVUGOvKC+uiWDCHoicjNZsTQu9mwG1JtSJh7khV7FjY5woJ8XY9ScGma62i5rnZpvTcq/uIXEw
Ec8sjciQWgCuAUT0Fp5GXuIWcRbVXc2mI8TO0y/jY2phtjbOj9/RUbLYp0hTLxxsSYHPpi0sQXpl
HXPibsSkRoIkMg5IAC5meQk2ree4mqWbT5rA3O6upeb3ylbgyDMgVY0Ln9ZWU/eqPePMxY8eykG7
5K6/ukCo1G9MzWRic+RXP/u//oKp7AkJ4y/keoZm3kxTNktQzFUXe8q3vMbUGbqWEt0WXGtxBF//
aL+7FyuAUMzDSvh9N9dkkjOLnisxDdzAuUgD1Ol8HVRbsfhlSycr2Kq4XK5TzoICq4VpLDyb8QJn
3NvafgjGgsvs1DB5kaCMMXV1o+Axkyhxy9kMp3VWOiS7wHqrHFXHl9cQDLfpM8tDv4AIR78/8guq
YY+wQ5b/6iCtEVZ/gOTvIVoQCMWsD3B5Pt2lvZWcZAcK/pY4S6z/Fwlj1vOoITwrY6aT4yuXzF5Y
/elMBN3L+1/lwESpu0TfnpxIARAwTUp5ARBnVIwBsSI7+VlEd5itTjCkZ/2Cmzdgwu/WHh3M+jDB
0Aa6YKmbNWTnqmb/c1VTbsB1WsVb4x0pD0H9/WJELHodTfMWzgVq02asAptSm1kDUncVfq85VVvV
IltmE8XNHSYLT80PH7AT3Fjt5+xAbicQVqtv6TW0A1vNpcigc6SPU2PKVt2L/3a5vnDd3DVKsZyA
hpEUNlnw3xAogo7EpdMcSaDLmJKgEnD0XbxDcvWmTbDgDAz3f31FUKy7eSdEIzaVF4uE91hpoq2I
eFuNX9n9SrouMWiaFMUsvfMz7+vHfdfhU6zt+Whl6Ma3/S5a91NSH1myS9wfoHi1Wh55ai4QQ+9U
UOmWBie1/bHb4Fk/ai2mYaXBQgYGn+9Wv06d+g2dKJOXsToYeVD5DHXvkh0uJucEtQRZ3wTTZyp3
j4m3CD2XG/QbK3zK7sw0ZKxLAvejeA77hXqMrAosZ3rHQNMFoe0E7SGPwn3St9cAljVIqqKNw2Tj
NVvaforb3uqSZYqINIKaJ0S9gB9TYsmmCh/FjYVTTrDXsDVh09zq0VxioyRmEXDLD3J3yASeRl91
MVpVfAnEkaJN+fhMCoBJLmXdiGYsBxnE35gDqQjrNlA6WN2aZwe4vsg6vHpSOE0+zROqMdjjyuj0
1dGT+wd1VRRH6+XHcCumeJCErnImqN66DpBpxx6/7Msf8oSSKJQOgSAmnUriBlrLE3FTtnbfHbVn
I38hoRnkp9jVugTDoiz6xWRa4M4NNW47YTz0HciDlXI89eVV71lZM9D4yyYGnEuy0qezhULj1bcF
dJ7qHkN8ZA0IXpetug6VyBL7yBBKagmQ1DE3uKkl+evsTe1b06Ib2YWPDWpjXcmgaHp6hsSve2T/
ACyGalD9Rlyss8EfhQgY+8l++uTbodCeNXc17abiR8ON8tTcrkqNF5z/A+dahnAkbZawRa+c6abl
JfQL+i6MJBWf/HE0/WOLa0QVoKU6/PnDzwgjenNyKqATj0OC520JpD3vqi+MXzId42oExtolMPw7
klMSTJAugm1IFMaayb63qnJDOWaCYg0cOOK6/UlW8lgkldJDJX9oxhYIp0bzomLAummpq4/aL/cL
qfI61RSUp3wLk73DZTRwfkg6bMz0jRvxteLIWizyNaqvzmRHvDdiPu3GapqQKyWzj+QoDnX38wIJ
9Uv5VIXd+POMxuF9cH8o+Rcck/idrTUD0+sAimnBFTq94dEkvplVt+EkObd8yV8xoRHRqFzfjmmq
+e1DP3UK7XchPL2YKN+QOjZUWWsIIBYUn379B0RoF10kENqDrYpQDe0c/Zi7YjPgGVDgg1Bu3hbd
DxfXoUlQYBKQQgSGIJzgz/S3GeH6kNTnmyihH/mXIDI62E5mFTZf7ExRcKW4bm5HwmzbqtPSQeqv
b16v6m/CUl4xU7o3a9pz6dAKEf8tculjgPxtkW3VCdrjwceib0GWshJGdW7UjTprlQwXydNU8ILt
+Jzdpht05PrDabecEkcvhlCCVuIK5ydugej6ad6F3sqg5xzSazp7L/SoUOGaVWnN3NOiuNSYEwEs
ziHPHa3ArDx/GEFrB7ZiuaN6v3rMm3PVm3GgGbAdcWqLEpu5z3paF9y+Jv9GV47xx6m5M2CDHs5A
Z7EPo/oJa4CXo6ivegnWOAsZV/07QotPixoJHrokm7pT3CI20XeXE52WVHLCCMDvDCsMCJbFaKF9
fDsHVi0Ev4pSNqADclEVeDtFuq0C0Trk0L03bxR+TAeRY33JWOkfPrDfkMftOrQyvIbgN5FhwX5D
VLwzvLnfs4gnpnRx+PbV//fxtMMjItbyMcFJt+rG+PO4+t51CJBHlMgoFK+w9ClPQjmjQcp5nb/+
HCnQ4OwQZkKTeg5GPt8GCzay9GYgpummFeE64tzOvAVS40dH90n+cD0sdqIC4qvQlRUE5T4nvfBq
l7bpP7rrh7XHTuyK3CHxxKkLH8NPywU/uvzsWmOuNpHjE2BjVUPi6uvBuFIngrUVNiQDn1f4PfJh
StQHR0xRK+VOS1I4Zxk2wAwW8XFtIDQtZO9zbQ6LfW8KNrEYmwN2ypnnTz4yHb+45b8ER8abmGZ3
aRfpVuoRQA1hk4+NNKl36rZzhFhj/FEFENcux14xu36DEGJc9vikxztR1202Kxrc32fgJGNnNm4/
mZpTSR2SdRZkmrqoYDce/E7lg3MzSKBbg+Mp8Oq3EYOQ4+mWtzNUB2Vb813iZdLGTKwON4iRY8bS
ow/Tr0hohRxESx/oMcx2xoJqONFogKAApFo9sGl4QtZxVf5Lu8TvnLqvYPNbdGAdrJU4BJK7clqW
Qk+gV8dK6Vt3EpVpZk7hKN/8YhOxLyiqmHds33IjFN2XM7ahF8ZU4yEQbzim+RJxj22MBvqzrpMs
I6RUHLcrsBX0ll7AgKIyxwm4kiySDMZSPG5klqVqFzucjKKhRbscH1KOG4ZiMM6kLpAX70G97Yig
tiyVbsQ2tBpKP+Yqnmy2PFa1SMfKfS0kuplFVZMwhc5riGDA4BkR2+7XW2xS2j985hzo34qXqzqV
Vp1/k2LLbqVkKAgWY5nqG1hfwXiePgJPQ+mIcjK5lYenN8NvvCbgsE1R1p7ykxWsIqImq5/BWYai
kc05dyeUXGEHEbjKYm/BFf8pRJrFt46dBbF6vsudyryCGCZTS8lzPkzm/kPqqKgyD0/4L5emi2Si
LdBlmhdTord9qNi5062vkrVAqX5brEaxkq30g8hviORP2ieILOECU6AAZuEhuU6nBZWFWll1JHrD
2OjGtjt+AqIMqxtwx/n9gJZwjhG8AG8k8sIqqX4haRUu74ndiqfkokSZMhuuA9N8FND1MAp4jNVk
wLXqday9KW24NfqVFfV2kc8h6vnDGIq9xXqkaVBU6HF0HrXxUJEr+OofpXmYQsLqKFxySVH1p1W3
l7nIb+41cePBV19MqOLBg6PplwbGfesLhFs4JT4DwosNJw82wB/0KhQ+jA8Z+wYYwQIbITAQ57Ow
0tgoRsmS67vyq1QpfSpbRAWaMHCFF35mxi9lQTgGJ4wATl3n0vlcy2nRMwm5fOAWBtvEMSLKBQSL
a8/zJVTVBDwEHU7kILb1Kd3suh/1sXGMUosTT9UEVzFXmRMumRu2pERT9S3cg+SrGCIT+7EIgbyW
LikXYt0efknmMiHy051K4+ciXSS8/j52Us7LxjnuY2rnJ80emCQaKt3sbB2JTGymp4zU/dGLEEjT
tukAaEbZfNjjZBW3FZlOqI4Y7ojrB/rc/HBWias32erIKZovlVf5qRvpWtoYdg/WXYvZPTbbegqV
SpcT2ncxlD00BbwDFXmYs8tHzm95exg47l3XSGYIl064CwXYO2t0ICrW84qIUD844spojShPdRAg
7INJkjotzceDI8mfo60WTryuwms8h+AVQ6FWBd/ZoSfVkhOJJI1aaO/vRCzr1EvuFYkVgveGNiW3
Hiug4YFpCn6oduzaVt5sykts63wldimrPWlMkEyd8XZIO8xiZX35o+UJm8r5w2ZKT6glB5fIKR4G
2h5LcPI89SmtZOAvrDDb5a9fRCwwbhGX1L8/sVGLa/oPccUjtJtOlgHXg3BoYZ0iBgkD1dhJxWrm
L1eReNKXMdWfeqFrQviAyZb5h9135qRiPqTCvhsSL8c7D93AFgWFm5B8hb8HD3FobWx3EvIQMCd7
OPuU5AwAr+0exur10RhSbYviXRILoFJVEGIpXTap9q8VOjQ1542N9nR02C+cQLqUGrTwNK2KApKf
4/bvD6Hdu+cXbUP678ScXretyY4C9znC80TQ4Wu8bsuaSuxfIt/3olC8aw4eaN1OcWbo5x1oU56K
JSuNEL2VI0sZHtFkQcA0UXd4eI4+VZD3v0Vwj6oXRdOyiOVrQVlN3weiHVr2iK+++b7Xn1MtNM7C
CEuAbAyPhcVl+9DOmAhvnNUFtvo2GIsc8ibf5aLyam5BqbqyQOFW7bfWZZYzDpzPRWNz4MhczrHT
UixWmpVLod+OhHVVBXTNkLpTNknYWP8f7FDvJO8YS7Bugm4BJoc8/2etGG/IxMnPE2XM5XP/FC1T
SGh5qyAVFUP0c6uWQza8i+jrYJHRBZkjcV5ep/8byHGKCUCkHy2m0DVY/Y6N16u6ket/NQBW6G3j
Ykj72cWbkGUGfAtFeFJ/Rk174s6fdxukeISiXPCXX0u9nqbqy3xPSi9qQFiEBrjp6KRF0noWEVSg
mWHv+mnazWIfFGu0BUjWZ4Rib5LBZllSmt0UjYCpbH0K3lEXJQlAPigtULEMRSJYx8evcDphb5QL
fhHvZr8eqEl8xY//sSSiPTSKI5VqjRGU8x1WxOyYGZx1mQKwWzmqYDYasd8F7vBwolahlW1ME1mC
v7ZswDP3QlkyfwYnq9qPXaHBbLoLIOQuNWhKrVyO1C3KpAsS3tYXXDSy1ryqBwCv+/6OwMR6jcDe
xGPRntoo1zlEWoRWbFwzBGJdaS3rfNBk7+CvP/3BESiLSavdxWagSWaOEd4zxaS4AC+hdz69uvUu
syovJVFZoOO8PZ31AL6WE/p9pvbCVHSVsXKDPuQy8hrZSVCxSlinrpFdvycZkKc/olxMR+fEw0im
khNUgeCnGM5YHjytqamDxIlVI67HUqH8ATtstBEKcS0npSaYvkBdIhe5z71aaDB0GfzWMlRqp3+i
8sPAymGiOqurN/ailda5GNJP67bdMXP1nE4EKbH5z1JfOD5R+/16ni5f4FzSs+J4wKxbV0XlBdaP
bopv7FeIlzSTxhEiVaVH7CftRzPAUArRCcve6AXvQtA8856RAW/M7AEj/IMK66/Cp7OKHvPlpJaF
PGK//nrXpMD1UrEtRSdvOCBNab3XJxX4MPdAnX3taR4NbQVSrXaXX9xsz7L2zxVn01iLewoOXJh2
cvPS5BqMbfRxAttflmUYvCfuMKaEube3votPujKT7JF3vVv6C8RNWQR3nw3gbOSTz9CWlTDlstMv
VpCjzKcNn39ceZXGjZWgJI2kkyZFCH2K9oPO7XmJygokNXbLMRuZpW/ZwgNDChh40AFP6qG/2rUD
kX4FAsdY2xUQhW28RtHgZ839qdZIY1jsPqvfK2VhaL4+gb5Gx7Y2pgAtpvRTYIVYz4CgPIEMHakA
wVgITjVS5nnqk86sXtvQdhJHGrmaCQHFjwHqFEMQgI94+ZhLF3st/LQDD9r9AZ8Y+CZDUWKO9yiN
d347w5SzLumaigAvhPPMeT3A4vcxxB0nN91oxoqoA3/Cbaya38JYwHOtZcRzicg2Ixe6nAzMC6GQ
HkitEY2F2XdJlZo1lk1U5r4HIM2JYwBk4CGKaguqlqHkFb0W4kjbGh2vRBTbC6dbbtz9wTF9fnFT
uNy8gJV5PNfJ/SUDDgbpiyRjbqgUD0iPWr9d97DmArm10Nb0wsZv7MWQhsWsSVD2I99yy3Hst28C
f27CevbXfpV+mi7sLzUt6LsU36Oig+lOyQsui1wxW8sec62GiA7OANETG3D2qkrsDDXe/ypxKl6J
M2WWM+7dRJj0NtwDPMDcydJk6rVm0m86bQwbjlKEVEpmUbzYlIwdjBzaOZq4+MGPbuno3s6CyGX4
DXezn0Hk78kF83vz2xG1bydFhX8RLP0+xf0JRpkto+XCH0696wredWLq42+JqvJTOyK1ESr5ZfJM
bRpNoqc9Xi53oYellhgNzh9Ja/+wW7+fyOL6cCYfPyzwtbpPlnnTnZ0CP93Z4nmPTu2+muVjI8Hn
s4D3LVukLKiGKq/c6vtONqND1ZZ7Jkep6T5gBv41s4W5dOxlwpl+AZHv5ziQr5baAez2jWCgu48m
lW2/w5kYqX2Jb2pnoAFIAHMRP9imLwDYAocCGW6OHbB+qQpeDyi+Fiz1P76g4xKNTHU5QjXB8V+X
xpN1iaY7UvAo3uLw6jEGQEFkH2YtY748D00HX8inRBWw7SBjH6wPMRFG2KS6B9WYrvNC/lWNMbp3
agMN4SiRPP03gXsPt2/vIKDJphF1c/O3+2AJyVZTrjNTXMUEPJyzno6fYMCSFHurfZxPLP4UxQFy
ZoKNUOTbaLZfLdqoAJBwf23bpPUbPcXZuPhEdyqjHvuG6C3Luh3brDU8CTSwxP3N5we1A1XQCgb3
RFl7/g7+qNqL3hZb5MUFIWPjLLJtANvyYMWZAl3YXPgD3mMzR97N0PHgM2HCyUjts3z/ZmXXUSjW
OZaSbwbrBLcVNuqPJ7NO5cTUD6jX/WXvq48UZU7StmNdAAEaVOkOquXay2dFGHneh9mWRIjBgM0c
S1BpsoQqRNyUGu9cj5/Jnn6X6yrN7VVjFTfghQjBhptpm4VXbwKmkfGcJ8Wr3dtgq6g/uRVNwPPl
5r3hAHzWOox9j4M3GRmTZcdfdAZcjoHOQjvBRozrA/kHBqGmaOIEmtLafH8cqs6Wv7i8prbNHUvz
CwG3SAz1RILyFMJPfL81ECiIHIBXpaVzJtWgd9+cyDsPgCR7WwA1+wQqcZnU1JTwO0rDN9kIhX0O
ey8yEpFoGaUL3CRhc9Rd7mKN4NOzDMCDczilAa9G2MBuU6z4Ekf2I+ZJVTRzgByZ/JXxNRKLRPSZ
RaSlJ7iRwOAdi+e6cKvfgN+21haKLH1XA2G8Nu9FHdxKFsOSGJAcpSxD3mpREWFHfZXr9MFBQfnc
OubyaHhEy6HswH52FlBR8xTsvu1brVoQcO6/1DAy8J4+6wgB/MCbT/Gm0Nub68UNAiq7zZ5vXYPg
n3HuUaGpml/9PbP9kPrRZjZ2f95P5OJvbFwvc+0po5JqFFyT7jxK5Qkz+cDVJZWCHF6vrlDrW5fL
QbJNe7gXIOS5HsCg7XKBcCPqCAY1D0hwRk9HF2PuK0I4U63k3CiMgJ0bayIr6earZbXWnJf0AUeo
GsNGeHAqYaic+GoY5yBvIMCJYFlK7sdbPWhHoLyDHW98Ky2qxWkOYwo7Zrt/atmPihJM9PtXpkBn
UvWaDg+ha+CLMjoBuOqEB4SsQ+V00fevRIYcieSpVwPc1/zBqdiVkEnsQsCx+4doASEFqz0QaOw1
MUSg9WreemECFd5tNtKqIIOpmt50KEaBn4AmXuEloHtCAOpCnHme+ndnm0tZJ+6MoyKTja8LDfXz
9acMhh7NudpMQV1EgE6XgKs5yUwAcwVHcZUk7lmaevGP+y+RT7iT083ku71h/XsN4qMufJsSKKnl
lUcyEfxZ0tioTPcnGpTfRMarVmcVX9nOsEvgMnhGUKoazsUsbGVnMTC+4QLw1g6UyeV24g3x/dLn
AFCjyRkpje+7Vp0qQzEp4EXPK8nJPpmmLVYG6vSi0bpMLKeXGMhHW9XZJyDFI9CtOozoMzRBBka8
7meROaiMCk3NK/6FrPbK9XPW5JU7al+0H1Dmwqkuvn089NgltbWZ28WgzixXzNcvr4CeUBTzEOgu
i7i+Zqk5YF83VO/Fg7xBaMlg+q8Akh+7js017Y1ccfk+h9WQgZkyYWmcYrtAG2fORLuX7SebANmc
BsrGYruav3gXQ2zgcxIKCS5RH8dTmXX6QbmFDN3bG7JMBxXkv+x8didFMJ9j18H53kZdTO7BIA4b
9cgrGTIfZteboDk5JctBsjvkT8hcrRBQoJnkHO4S4T9r2UqRKKgzHpXXe698GoZIaNIlpjcTA6tp
1iMEQPr2UgFrKFjlfPf+v1C5nA226/LY1oRIPZrifxTf9hevVbSNx6QYW+qBBegDGDumQIBk05j5
/ETQLUVEaeoNkkyGAxzb2ScOQ0qjSbhj96SQ7ZE7ohtll5fNT9nvSGnA+USJzYViBOlAzyq6/xIR
hUkoPsiATPqAJD+6y3/KlF/5WCc55xGoBXbxuFFk310isAhPCowxYMpIUCrYPYv4bml4WZ7z0IAx
R9ci6B8Hl6q5UwfTHcLA7NNmzDxM0R8fnp+T86vikIYrH73TTKzvdXRtNSBkemb4qNrX6tcuxI2e
dZT9f1UHsTEAixQCKncCBjFk0dVkmeK1817jMDeRYPPXr9vOKxtpCxCA8uTGygGw46vyhVSLs0e4
FNSVAYoIMf6wFIgdos7PsExLXaVwJ22Q9SDrL2UqCzI//ArA0piwhxl+uapxZf9RspSfzej/WOoG
ksKax/F04jGhUFF9Px5sLIo/oPY2FHxZ0ctkVlGEtaqOuwyppzPLmIQI/+3TTX3Etst9CnRKHYki
VGp8Se7yNhp8lpmraRcXgwrABcS8riHCnaR/7XPvBfashBc0WGg6diKJPDcpJ05aNe7PBYlGimqD
j/xbT/gmq4yypn8beNIhgtzAe4BD00SKH0XkA3yDfQV47WrSe4jWN4woghh34csxebJGkQ3xrqeZ
SM2bjgg29QOj1kJvtPNuLktYPSVXFYjIqVs062fbStzVGO7lGyjkoZbUbX8cj3Sy+NQCD+g8eE6o
ZP2z39WIWx0pksz1vDGUsueAmPKaZdOU0mxOzuelDfqLJTEl7uEMohU5PgB+qLicIH6DVc2GJo3N
h0MwbWN7S7DVt3bjvOghUq91gE1GHcaMgAzi7gTe59Z+TT88adCGIR8uZO7uyocUzrlm7DX73yf4
3XbcvguqoQENQqC+DxPLSqCIvwnaNnUjX1d7c13EoN6xRAsqrW08yx2vB/PEWfFp/CreqiDSf2BJ
9HiD+TX7sjHyjhRfW4HEWDTYJh5hf0XCLK/sc3e5GN1kEPGbzJObFplVtQoxhykCcod6WduQv72L
lBaO+GUYTgoKJwpGGHMypwdcJoKu8BThyEW+kfhjMXuLiIGhNc1d/NLoxfZNyMj0D0OY9p7zytQn
Fsd3I+/uu7mAcZ47t+kh/EMvUquajIQcNhivDAbsaTWDKg0hMUDubKe0TzKMiKiu+XzfjhR/qq2Y
rUDZXjnwTHTMS5/Kmfi0tXQfSUXLNU1/CnMhTxQvt+IOmBYdDuiKcoLpF+HWzag/KgeFkAFYCdi6
eoK78/kT/DCMW1r7IKUotx6K4xaIFnOplXEmUW9lKgSXMPCUqd/YnX+ghmfc2FbtwLs3gE+J5dTP
RuXjNnCS3uifIQqHiuxqUaiCMjAZsnE4uxAbf5hw1DSOehu+ZgGxubQnSHcRP95BxndakduBNhyS
uXZKtctSdVSo24rgwtu8VN8U1gUF9yuybdc1USaDp/lbwBsgnoh/oDl7X4s2/p2L2Tqd5iFclWqN
BUuBVDfrtofVhrl2vnKDtOEgGsHAPlDERWCuIshSdZVRImivr7mUU7qnsExoCxYDuK4E8vKayQwr
2FtForJSDjlJF6NlBvtzCLc0weLc2zzZH9LD2S9XeOX8lnRCWdN7WluOAz6Rf0oiMCM/njOInXqw
9HvJlX2y1x7C0fNCPU4O/O0omv0lRHvkobHksmrxi1PYJ540PIMIuC+w7fweCVUlxq+NQqOYZiuc
1jdPR0ppTBMvkEhd/PJbIMQLC69rbdPeAuqXCwsJE1njxbq3sQC2TdCfHv1wT6z7Vmg2/+6+caAr
qkqPkAJU5LV3HO2NyyG5n40ucs/zsXS3bhZKdTAfbBVac5rr9AEGDc/4EHuWKYsZu7Ewd/ag5E03
pDgyHes41Ekb2RqTeovQQfzbVaYweFBpW4tWBvG+aKjZk5M+XSdVUr2utc+rYG1xDy8EMe2NOOTI
sNNiPb1RZFKvbbDAExw2V9tLz6mtzMJ4+TcxdV89ghik0r8Zd95NF6knCKw9E4S4a21NPJt9u8Sl
574/IWiZ5hLN9+iqpIGVoszvb62UJvHbCVe6aZRyMP/1Bv/US+HOoE32SD0iSnnr0metl49bYsNZ
GbdTF8wr3U7Y1VwOAy/HGbOHpJxHg+BwSY5nVg0tx6G+CTxWLmlpu1UBPbtOF830Qc0HjmrvBEaK
G/hzSjRQIzNatSM1Ow8z+b8tiazReKRTgXnKCqNuub2Ej2DU/x1QNWwk8vkk5RCjcsaXqIjVcnFU
tOzFTynzcplK4YdFAplbzsm2XATUNsyRjG+VBMTZANutl2XuD/tdrI5skpwK5JfilAFgQWdTwGqK
2gTSBvb3JYy6Nl24rJzT/j/wdizgtATlW5IoNTcz1M2EEyWx/OoZ2ugRJuikOdRGf8ZARhIRj93Q
2uC2s0Ma5SdurfShprCxg57wDZsRUEst+jG64uyUcfppwD+TWsO1OUi5UvT+/DJBbDsC9lygHjWG
43HSvoOdXENsG2kPwfbKqN+nWf2MF5hgGKAZtIiygSrlHEArl5EcbMgUKPv+yGzo0S75PDpvL7Dn
BAPLBYeCvFyD1h+RfySnzCSIrhKrI8hDdjzOrdyEykuE9gNkFBy2UH6F9PBQBUdjee+d4MDc2pzY
i5pNQX9bOjwCI22SNzSzdUgSvBKUz0Na062x5hDKurKUhgYd+5b0DLWwo25eDl0okfQTMyPlTTY+
ekQlTfyUfvBuydCKe6j1hXLnf3ubwrtN3dLbBubgMgXT8DyHAuQm44KFJOdhO8eubqhixSaVxsKG
buGiv9Azs7E8RRMGhMmA7QRiaW1sOvVsfESau4mO5A0NfDPJV+b7lUGs7mPuUd9q+v5SlFENvUwE
LmNIxcRsnIXDk9hTiZfpqDTn/ClDpS48sY+gnY8hjy34BdL/2Wmi5E2S6joOv53Wh3BZay/LygAS
90raZQ710KyZB84n6zkz9lUIM+tZqkVnTbS4XD62PqkM6DzQaCR7w7Ctydw6bR0C4jeHod0MTADa
5/cgLL3zUJcSJ1+YyScLfWa8BBPud0M2XiaPL6wtlNFkufFbGurWAkHgHL4FBrbRZYeBcHTLT3mU
TJcCYEoxlr7GAtKJl9pOeWBRdwniARn+Aj33AC3b3j3O9a+31FZByHVXFkWoiz/ntfRq2ZQhSMLN
656hBxS6GF1UO66A2MOALxuBtN60pYO7vTaMuD+zxgc1Oac/lU+PBMhOupjuLNQnm0FO+fX8wxTT
RBNDr9gpPSRg/0Pq6N/ZWrjIwc5MOVF+QveB91YmkgAabyn1QrF/XtvRReXq1tC5M33dwFkkcnef
W20EkeBA+KLBN/lqMLPfaTz8QWx9Llq0XnNiLBUt2vv9GGVePvrMuyFQAybZltGm4twdiQYeXfz5
oFe3UhBxqp+UPy6IMprzSdpEWpL5oFqy7oF/N6IA1qryTp9La/WXYPH/aksXlW5+MgVagBYdb7Qz
/bYELNk6yAwV0yqnUjTXvwoUFNqKDqHoj2jtAfYGhu5TYpG5PDR4bhAomznGCdKMiaq7Fqn0NvHB
4OAdBFZFXwvl1vdmUoX0fz/h04DXZb5sdnYCUpjAfg/walBAvmH+9VlZ0Lf8bammcbpw9i3E8sA7
hPNHKMWkOdc0iLS/m4r9LQxJfJRypkA6Ewdczk52h3U65/gtoAIxgRF4azsoIhKXmV8T9R/whHws
ER91oP1gz9IreTtlIQ+JpA2t/jVWdbZmfXFAilPOzUqZ5f2CRpL/LrmJvOXb5xn6gqIccsqW4mUD
kApv0tn8sPWz6Hy/laZWgbeiC0wWZYwB/f0rPrWYCGop4+GcXNda2NSDdI4dtrnxJ3QMigTAIcOD
+0Di3cyjh+tl1mTJhypHfeE4qL6ExNppezX3u7KFVLRnNu26lgLu/5QCSMOwZjeT9AS72e5757xb
oE/1sbizRO5h0KymA7WrQlnByiAmllcUcNVwqORK5IBsAu5hwd3vFTzY6kXf5nrlTXgfFGyfPu8t
+t8LIgvLDEXDEIjMx0rFwPuZk9eMk9sMg1Kf8/7dPguvCu7l63wLkcbEEM7I/EFn4opZVhTZJap7
E4JAgmubr8XyrB61drVQEot/lE/pPjNuY77Kc/nk8GwtTak9BadNotoHgOMJWjQP3xpiPoUDX1dB
evIioGIkqoPY9Wl2Ux1TvVqFOHA9uKZxlDr/CROcBlyDuXoPIp1/VzlLmutlTlJaEHwffQFJms33
uu0swmbNxtkduOorNTgtl2uOrHWtd212j+zAPejJM/W89et4Uv93RtelrS+ZM+i+4A4RE+Q6n1YZ
qrJ5AGWvfXCsJgyY1Mut8ibVbxYzMNOYlNXKS/rhiatotC9uM7kICj7c9GZUiNAFXa0mPMZ0xvop
mPwb33b1q/0BP3D3wX26HrNSdtluaWrBXiuvuEg3RjRFPM/YlKZDhubKwvHSkao9dFeQP0Ca3ydc
4HNO6A48JXUjgNcXbi60qA5dVD2TomgJNc/4KnI0Bmnuw7gGFg6lnY8Uh/1fqbNvs+ZAoWm6WU/Z
d3tR1KiayeSoxaugwenRXvQXS7MVwwpdxHMCPhoroNofnW+HA2LsA3V27vNwa+4tT3HaFGADvgVw
PztxMXVFTHHXna3z0/e8SOmUdIvs3qFrkotsZtwcRQvgLqSBij074j0FAyfUpRW053tvckAxvhFd
mSD8G5agCNbHQihQfy4VZes6x8kBkupTzsBBHpgFH/LMxKz0wUfTMmyPTLn42IsieOUzd09VQTpl
QSav1V2m5UOFZ6YsEoOz+SbaW+wLwvlJbRRfG6Ss7ou+qajQeaLsZFR/LcCL7qp9Y7SnPn19d+DI
0w4GderKZhnHY7CliVqGizZ+8lHK4VHR9pfkhCFwpGJOC/aGvdjjqOrGlwZ79KNfYKFZfLEdXV0G
ZGzyhQvl5kmFDRaWKcGDchlfeU+gEZ9r4brW2gm32U8iHIEeDSq09pwQBx8gVRNbBrMyANHzVw0Q
dBA0GQASihaaLLGoYtAnckrhCQd86/rjy5O0ghIbrRTxcmSm8hwV+r2xTDrUGi3EwcrVUx96qFJZ
ILnSPHW/r1w1vY6A+efpKqrG4e9h0uSfYyuPz9MfSvFY4x2xT8SRICGJZC+2sfrHRKFGmEiLUfdv
vBPF6xTBCNP0RRCDE6pRxXNPoeJv+SpFpEcYCtIWjY0VtS6TeasiXDSsf3txL6dA1bJ8/qr4sf89
f9Of/07p4wsgOya5kTXT4IsgZAB9X9uIgetRuE5NiEHLK5EcqdxhOAsw0uWoFZkvG6T+sYY0U+mj
Ug3/RhTodAfY7ZQrjcLTqG8WF/UlUTNnJMoLsa9dpZ9TdXVUS5evIfCvb9pF8+oy/3E+n5tTuY8E
c5C7BE/4n7riR4TyatJNVDi24d1wMRgk1JJKcmXqAJzFew5xNDn4IoM5vT90/Wjy5WpokfIvmYj+
3xxWx4dfdobD9eZ5iayMJgLpvt3BgTXvZT0OS9/VhXQAKJOlwEEaQyNWBNS5Dy/2hEggDTVx/qs/
keQnw62xuMXOIcg2aSj3mwrx00JfPf/jVpMpM++3Rhsv9I8ewewwed7LuZIh4lPONXYyUPbT/nQ6
gu2+BbiKY9Z8xS6tpoMVfpL62BymRiIhoURdDj9o/mhkn7VKRw3cSiEAiBvtu1sD4thMznpx44yZ
buz3ttCEY9UYupvayuPBljn2hGwEJyclnTaKGpcgfedV6Ai8uN3jhtq9PddSZ7iqEbSxbpYV4JDs
bxUVG/6N7rEinOJ4u2xPVp42osl36s2F94ee7TVnWJnx+9KjM61NBJ01lWyvQhVyzRr50TfvAwh2
m5cKkNDFO9fr8iWWiZwIuATuohTmzu/SfvX7GBbZi2Q7vbuZhOAGFlmEHqcU2YYWMR+FqVPVkLmI
zbJbSpCM+kgH8TDI9VQBwjeq/IUY9ImjYjbZFX09+NU89nSZyIZZuMjQr/90Y6sOt5ZDj2moScgC
9MthHvUx7VHSVzvHeCeQAyHn9qg4fNkJxF9mfbQhneIhmqNKwJvhpkO0ZlPhUn/0sgeocF3EhuQU
ojfdx4RkdH7KvXZ0wPFSZMh2PQKBvKkGXZz3VjZ0jJtvU2f//Z3Vvjdrvs4D/BDU2fXEqKlebIyK
O57pTUbvxbLgZu0a+7PL2+VOeqAD8BDZ+rd90xb9YdOW0Ft8+8N8s3ZuzqehwG0Bajgb+WmOpEsy
9g68j6o7OQP7WIXzXS0xrmWxUDdbH+swcfKgJThWNNqiY6tXBrNTxUzJ7NdxZkhxSHZj+oP9z+V6
3zziuy1p/Ozghweta3md6LGZClZPTiMtwqdsCfUBXa8NXPt/x7sjtOQFnBiu2+Jpbi8IsoK8eUlr
vRx2K8negR8GqpHREmKqKRhxtXiaeGf3N1sMrwTHVJlHBXkEB4QYq2hBkKSXy1ZQMau38AH5L7va
i8TpHzXc5EEl+hJ2ZjWN3zIIJMG5KL7y0hpynXoa6X3pj4c070+udvMvojs8B+fkFhs4Y4EeBi0E
XWF86RGC68hlmK032t6oPRYcYKTR1Ed1OhX0xAjsLJ9SAYeq1DY653IQ0k34f3/nzAzO4JaFxByF
7EU0xleOHPQifl6IjpFoz+6QehhU0yz+hvI2sURO9CrlCOO8y8zhC52qSMQ5cI6UwLoBe45QvfXU
+At2szzbx8cvS5L7G/LYqemNM1H+NZbY+j/lVGDzdXdab3rhvppJl/bM6oXgjquYuJyWVIClqVOC
e6l9X+3aCdl0z7rXL/N8sF/hKaEt4H5cxCoGUldwM8wETrTby6cH7hB2lrKGj/UtlSrJbNCCBRag
JXEv4cx/5thyGdkddkSMBhPmVfLfVGlNz8gfyRhqgHsvyf/hswqAyfNScodBO/qaks0dbeLyxTHs
pruhwCYFuJM7/BWufRXoGCce5XXP22Thn7r7DypjZoDaGwXWPVlr7sx0+oWlbA2HLNur/RQMo7P5
4BSnUaZkqanK2FDTsQl66me+JamFQXnckdIBxvb9yYkl/mqlt3XqlR3ZltFnSaM1q1nxEvPx0qrp
uzX0xPa7MKOpAZb0q0noOpaZnTaOUpqeHGrLzQ6lkR7ItM4rLYADXe+mFuK1vLxg1fIza1M4CH4A
qaH2micpH4dP4atKNkT9pv+Wb6/8BHS8ZK3Pdnu4P9RLE0DdfMXptNtw2X8xUNT4sYrtzzjLmU1/
xRwlC/OqLl1I4mGyM9YPeX4GxXDi6fJlAwKB/WOJjtsj3JQXBlssPQCpqe8N0rWivbRuE462NKOZ
wVCFIb12y/7ipQj3f5aRPuvPO3Ypjm2KZbdDQql9xgP+O63Rt2YY7MNpRAEUbtb/dv1CpXrFtL90
RPMxgWoA4h0xUzYGKpzaf6rqLHGw/VwCBmg2TwguUXlLWEeaDtwgvE+FZUdDBUVmzEJUpUEk98fh
erEFUrCLO0nSH8fUUw3ScNjx7TzD6q620g7YpBqMpRRHS4GOHxrW0orG6WuBy5xt2T0t/80EurLG
I5LyASp6lPIMj9eUNfXDkiBuPG8Oke9HCIhGaty83l++Ph/pswkc4f7foCsJx13cItvMHMQp1r3u
nubXWjtl9Yhal6JYPm+eG1lKcGvN3reQd64eR4iNPOSfUcEf6FQaELnzkHT15B4RhOqpB1BirLUc
aA2t71QWZNncZEsxiVfjDZIfcjM3TMpxdyNeGAMgKgcLE/Yp+ZEbkLrjCuK6xEn/s+KxT3lcLBnN
QvQ+hJeU4noFqnpHkvK/nhOncRf2WHjwNmQfbcKR89rqq9dmoTpmsoH0qhjq+n6yrA9ofFZBT40v
S9S9NhmOOKFb7Pr+6Xuq8WQxObx11/7hxBZv5kevE/SHWpY75aHrLNBG8kthVWifG6vGSLLQx+A9
mYtX4LxO8RjSWL1i1SyBxe1HBAs3gTRF8sUvdHtlrwwOd4ktUOuY4gPSO8lhZp/YQHmSzmbQARZg
sxuMcYrIsq+d1W76wmUeQoDYRjkV324lDUb4JspYECInikY0qv5AowoV4CEUIIgJg79QyEhHkvqY
IF3+QR2Q/mBphkRdo/i5nN3YlsIZjuJf7G3dNezvgheH8iJORAYciDkXcMBU7+uxgNIqusHfWnz6
O1eq+zRhZIDusEP5zP8Q8gZC7NxIlQY34CZfrqr2rXjFJpV+SC8oPv92W8jcDTRXcGiBCEPaRSI8
cbWRA84Fi0rfDYVSwpaJpBaVHUdII/VBoX4pIfPHwJ7GdaujcmJGmcSCe+MSnIL7K6gcKVkfskno
MOLi4MzIMGsCSHw2HmXZhBuI9WswFc7DW6GrdDtCGUhzQ0UqcYPPDHWSbDkBcNhcVLSBwPG/U3QT
cKeB68VDyTWM5zcIFwipTtUHxwj/SXGZeAJobGIuT/wdN1ebtXh3tICceyUPGMjvP6vQ4VvKTMLu
ftas56sI3RarkpRcbRROHUse5V6htDriwBV0AZSSGCvdlpxjPcNID2OLyyYfQWS/8cXvO5IXQft9
6BEEJpMS7ZcG1uIpKSuo+KVaJE8UUV+VoTpyYREozbWxaWgB/AYht1wKYLl7hdaoG7PMApP6vQXh
mVT2gTfjFHqgQ2MBWRrdmBLCsfd6j1uOAbPkhLhT/Vbju5AqWqE3XJKVZAhH4kAFUhmYQNQtOd57
vZyMN826VZa/uFmIPrJBIvhnGw1P0PklzzDb8FLiq5IAbowrIC3LbBJM8pc6HMu1VvI0HELqiC/h
GhOSm92+1UpRv1gczcVaORFtIMlXpLs5TIR+ehDHAPUSvvqYIn7BQBjluqiVxcb4bjZ5cqsCMRp7
9rAQZJuinIQzsXBcS3ewryo058c8ShI0rwBsHh6nL21u9NTjyR91l28SFWMQD8Nw7vlOy6EQTkcj
BdIyLhVY5m/B41ejcZb6jm+3PUtI8CqYPTo/OJdc/J/JjcoEK8GTggvYWl/xXywRyyaLm4XnxPRc
/zSZ1PzZwV5oJOhtSvm7TZSOgK8dUsIpkMgdZEz7IUwzwFkR4foLWozhUw0NeIT0//EVnjfahTcL
VgUNWcYH3vmblpN5tnjJ35xqn5VSyD4aR2TPCOv3wotkhiJ0JEdgoOv5j7f8hEJUlRaGSjd0HXNG
9kHxQEZINsKdcnPgiGN3k1hFkygGkB4a+7Xk7/SQ+MwZ+dtV+SZXqvkitKYSKPkkUisS8Vxj3Bpr
9sJnSuFL5B6cw0T67vLxdtiEznvssTObFW8ZYLHyPzP5IrY0DFooM34vqQ4k54VJb7UUp9Ozfd61
COfM2agOw0VaToW9u9wPI03Adt7S7P4g/zur447XSWd+GUXnlSnxFV40cYA/JwOBcOnkabQ79Uz4
rODrfI+JsdMj3onL0bgCpr3n2o+QAOSlG+rSnzRacZ3wlgTFrNvpT4dbd2D7DbPuxIGnHLALGH3w
jzJ4N2+90OBNnb1AfS6RIVIy5T/FIlBe+XtMimmazhSFrcmNpB8zgcS9pSUuzqww+JklopW4uLL8
fWz/A3JvI468Mj+9GdZJpP3d9fYOU+XNH9GZhPdvvBUXAVMUE8wtTmZx3XOwKA1H2je9grUBPkKx
B0s6SnmnZElZMgJ0nQZk18ll2viRvw/TZmT8QBJg/BPg8B/ZzoaeOk0OSxYckjNFHLM8X3c0ydUH
gzIN7O/kZosUFhXhtHfltEml1Pn/1Tspo/wG87o/UQEJV5x5MPFlF3+Pgna9+0iphsOd3pTTGw1I
uXihwKLeC2fEUQjlwOz7Jq1ZKitmYI+p/1VyVs8b3eAT3KbTYx6Dr4xoYSM7o96uE7cR8eDs/z5j
HD6WHzdszl9j0KKV+UaRgIHvJmyWsvo7zQ82LtOYYbH4nvOISE3bUtZqRv3CvR0VJsJy1DEyg1Vt
6qgFvttMOivOSps4BAHmYdhHbB5tB1z9z14d5olDH/F4iwiGxkoOno3W80OxyswlTLrYC1NNvtwE
MaLgG4aKwcwGOzhaYQJEwZeZtfRjf+o+D/SHd1Bx7XIG59JoT1M6mDQKzna29Q5XrpDQoLoq4ov6
UP4vKV33B7OnOOlkGMeO/scy7kdfP1gFcFkva/Ei527GDtr6maGRhUljDb5fo/L0yGToxOGHrBwv
1JybIx03uM2/UGl49mIu0+G8/fgrb9uP40YZlDUHagkljNNwgBcWsQ2eqhrGcCPHULUVEguO1lCM
ZocCw3lhGQ4HOka7fTqxtRCJYNY87iLXGt32s3MxFM5TNVN+2P8jOuP3AoC9AwPZ8nPshkwamJRD
P0CDeMZvxHDM1eMD3G7S53TCAs4+D6KEy0fD8qrxuXhX9LNTf7oqOgUChN+eq3bK/z0AjT4N4FDA
0JiUArUqCEY9MaKwQsDj06hIUu4MRp/pbDKvN4ZEfq2Rv84AIy4GOw0RChcPwCIu7EbCX03VZPRt
AHrHQ0SLEbwFCc2qGGRwhAKvLdZZzXgS7IIFlhhTljL0aR7Q847w/7LGJKShZ2ik/ACCV71TN9M1
/STQXnLI0hJ5CS3qlknqwfp0uoVJoFmyM07eXEYYLsSHHSJNgWRSDEQNVzgS8HfyuMVkIbnrwuw/
KWPICnukVrBWbv2ieMjPpVZays76QK6Z2guG7MYQOHAUM9yFAkU9CdXR95oCJ+CWUWY3UexWuOE2
zeJVjH1lszHgk5I3f3UDaICJqUeEqQ1ocZPkgU0C2stX+nujKOf39OrbuVniyTu2cpAPqCx0ReZC
BuRzy/Fs2+bw7QsU3ORvXD+DbH3HfOdkZ7IQ0IRzxYVarmTpwJTUbqNLaLs5u7EQF8IOuGpiGINe
zSuEMJl6MzMnuAHscWsYQzzo1ODn5PnBJVnV8CNQ13qEZssjIRAQ645e2zZvQ3MqeE7lg8Ko38+x
UkrmLSLKbvJhGqfc8ctNbgQi5XdZs8VKe0vwPqMmHYh89L8HXF3nRiTf4JmCEJ3dF1+XcBmV847W
16apMIv/E6dbgczfZQjv6awjSe2/gKn3G0fNzhXYGxfgDgFV/978qWw1/u4F/a9vgUBAGIIhMwqu
Qql/5B9RoexX88pCY2yEfECT1A8EsIC6CUjU10pkvqy6Sjc7eFED+SCutpBOxA61reau+qcWEE5c
rrlxmxLISKAf67MISpez5daZhPJQU4iNkuwn16Bg7g8hEbiDJN91a/aZ3okcztYfkHvkNMcLD1VY
7iS6142BmCKusIM/6QYhEoMuTzRduVe+NHI3FMgaSawhc2SrPKFVLH0UYBxU5b1PZGxVMuhSwaY8
3502EGNAoCDZ5povzmzSzb4CzD3hnVJFPduaIrwQ+VMdqsXxQ4x+vRXRlYrnPp9vbvZxSJ5icqAG
LTSRRg9PVaQgh8t6XKSoS3IhYS3RnGaiw6ke2iS2Ma9Bk6FJYYJdisvWxJKCBEzED0miwAR25f/s
jcWSJGcVRjcAhfVqsQQvtctq5Urj3iN+/0SfvGvaqgH8GnAzanVYu8cjg1zyQRj9Vvsj7y58PFwv
ORPI0m1Gt97hnlSn/n50ngc979w7YDB+z9ojVFvr1RPUJATqCiHofCI5XRolrNzCK66tfVPui3+S
0HozqlXLi2nlX5B0Wqo0R6YEGoATcN8GuQVBp/qRbx6qxLlMZVedJA6SZSfBk5uYMXBpfhzvzhUm
Oms/RPi0LvQpykxSeDTg3H+9qgN5tu2zs5a6Dvn8lI9eprfMSws3N7oumCYXiPbTF92tP0sxYxGa
D/geefd/MmDGR39/E2pzh68lDlR4ihPSidKvAKsCep3JTY9KrdYLo6ywPXAYREIfdKw2anuLiYMu
EM2KOH/KgPo7KVKr0Jy1j4VEgBvVaDd4fqJAamlNzB8ZCqIW9I9I7fG0xvkZCZG/pZ0xX6XMydlw
o8oUmtxk88rsLTk6Of31MT4MuO0Ddy8I08kweACfI6V3r3giRTzjYTE55nkgfRiXELjZIuizytOh
4DfxchegzeSvPs62MMxB/0KxhQFGDF1ZPz+0oo666gsqu5HokEGhvqHEixjUnNSxL+q7hy1BTdWc
jZC2PoEz6zwy+ZsskW0U2F/RPh6vkTsjiwqBvVO3lkzzPtG0HT2hfbQkZ+OGMFfQ9zvxGzwgvmoS
eOVlkNtx/u/TGkQILbbeNM4OK2+OZqFubwn0iVtCqQCJjyceSib+SXPnpwsqrrDxtYGUn0uAX+HC
3sFn23x1ju9FNbUuvUiv+BL5bRetvspCcpzsP0yM3SJekzli2E0v7TnlxPLfVurP/vlyAN1aPHQU
vtmVhdLzmZybxEAnQdE9F/zvfl7lGvg3m9ndx9P6sN6mSbdlf8LITJsvpQWgxIvec4VlU2wxKp2F
CHxxFC9i0QVJ4QSsfvVb0463Nyji/CpHx+UhLK0C7ve2atDnPkaoWWblaISKCYEuju3b4YHL/dhH
ABKr4oPJif2ed7YmMt8jfTr4yzn67QaW7Wx/avc5kMb5B5r2aE+JrhB9LuEovK6qEjf5ukaRGavv
NhqdrmhqvKDfW5rjyc7xhsszlv23EkdNnm63+B8R9qlDgEc2pPk68P8Vn2gdcVhHTrilKjxMCPrw
96ym3uRNR3c5Xv+kU6K79niHJGCpuwPl9dCNKouuAsAB1t8+ToOVfibFqtFxbkRYmqa6v9xfTjla
cUEZ2CpcI3ySPOy5dUUQLT6eHqYcg49FiXxqPj/9b5rkUs1f4mH5I0LPuuYL0/ic+O4YnIQr4GPn
UpgPUznS8yu6qKxNuSkoIRgGeheH24XBz1fZt7B99Lr0wUKfbTh+P6Ihtw9k4xdUWwoUyJKHTekD
DHbSC6dPlywHJKv4OUezAgKBVjRkm0/kLfMSLJ3PAhN18YZkqdHpiqHr6hUx3HdIyIpqrKyhsnw6
to3PcMEYnIqgFYq+SwTImhIiWLOwv39q332XtqCylBC3oXaN09bTdMIOQHVctVgBGvPazyqH2BYy
6AqAb0swD5sppv3635rGOyUj1EDnVH8zaUlR/CICSKM1tiq1cCP1vF+r8ctq+DfYYGcaiVnuV4y1
sYBeL6myVN4aPTwz5dGd4libiJIYvdB4XFovthq59yYLITo+Uej6kQ0VNZQWADqfkQzrd+wALYa3
pS0JykNO+lVTbtYE6jCjTXeD/ySucVpG8vfNwMDwh48aRnGh1qYk1usDBABqlt/4aeJWk4f9Iqxc
YUDVPiYMoDwDrR/mIASYEZmK+Qt2r7ppIvjraro7NYkyFHby3dGGFog3jEtpIHOAqMSejFcLUtv/
f56UbujQYL/0vKv9bsIHPlV/bPUBetcnFeU+f6auGCqkaXMFG7uNDmoEOKq36tT6pasicKp30ChN
TLfEvZr89pQbEN2DGIScw6CQngnEhTU31buM9UNjDQXdjwIJPb8DwX8MeEUUJxz3r30d3MFDvsWJ
wLi78xmyvoIg00PyZ6g8wRlI/LYUJrdQK7pBZh4ZdJ4Ru5SCGvaELUjacQ+Eaos0x6tXCe7tLgzS
2nNJgiWFsaTqwom/BaUYjDAntOXavuXTu3CxAwCfSP9grYqPWCNjY+NnvEE3ltnySlv2lXX+GFL/
525dcrga4MdZM8M8Nzf2VSgBriNfe6AEwxbz0OJ+obl5km14Rd1pOeqV121qAuPaNoAbbDnMImFg
JA5nQ36KcZq4I+7HTazxCPKpsOnxLie5kepIzi7VA7l5p4Kr/gBNZZ0f5cn+z4GIFF2u8oy6pcfO
BVsbq2sajnCh9gnWpt/+PwDTMJSVrU8Zw0QInLxaVXlQ6aJ6wa7s8rXOMAsMP8sE6rlsSIvwS/X0
pGKQFNpcgn494xzH9yFgenmE9PJi4IRp5Fet6pTAT49ZxrSML51dR2TJYcOz8y6juUVdyG2LD5iy
vEc8cZJubWaW96iVDtWFzO/zfQWxF8q9ee7Jq1Lm2gk=
`pragma protect end_protected
