// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rTezKRheAwQQF9et/YDSNQ+qcpKbxaRSnEhI3PnSpe0StaF1fMPfO78MN40N0fA5
Y6O3F7VxJDt+o5Rix85XslP1UlGM/CGN/bh0RWX/JpCcRJhu3/Zgg+qpYS0D33Kb
gulYH3TGqVu2/AQUV6MUteEX1UAno53lWtKlLG6uIJI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7280)
t3bjeaae6QO8Y0APqdLCVyvGMJeiZmCzA00hAcFTF4fPBqqdAemNBA2bSu8sBscT
KjpTtzmYVA4Dub0Wc2/NQ4OU4/fP90yif44LpyIoQP29vgLYQSTx1+AFHmr+Xu6g
tIkIdLCN5zhQyYNVauwpaYHu2rNe88bco95GLLtNi1TOiQNHvbcG5kkhRnNFStRb
5pv3c+Fjqod4NIYOOnDkRpYvmoyeF5tWFWVLMrqOp3f2kdirnJCZ2GlrtexyVwCp
7djblAA1lQr0bhKy7r+y6Z1KT//Z45OBtsFSU2VeDQm4UNKb1d41ASfJWEKNlRJb
L8MVHzLHTPW7ryZzZevzPO3OdnkdCjqF0B8DbkyCf1TcOlxqdegKCXKUu8+q7Bbl
LxeMbJh15/L/Z/gil9D8J3kmh6Vlj71/b6hEZlcYbQIDK4nFzeYYl36anJMQg+NX
ol+2GG5MsZsFpYP2/PIXszPj4HuXkpxjxYzLgwer5A8QNcxkHKpg+7bbq/+4XiT/
IBOvZlNFoQbDDU0BG9EYkWsZs5uQLzSRAk2bRPOyhrtvOl4QXmCU9zaePCi7t7Ol
EJWW/r8dt6Zr0XXOY/VPt5V7RjOp2ZPU9qKh3gllOYGPR1E0rJ9gnI2lw5RkKADs
AOR0yDQWpbWJ4UlNPGa14ZVblIrShwJJTWz3sc0In8nVk48tvIx71PGXqA+WXlGF
cOqhv8Ov6RBTR0Y8LbYOQFK+hoOea1CvOYx1hy1zZTu6Qwjt4iG4prcHcDt5mrSg
7XXmSc4L3qyBLmr0v7OLwz6G27Ac03iFbmJDbAdmSec8f19V1Cu8cnwi6aJ5Nt+t
Haycg7+VWfEmOf7i/6KAl+MzzhcQbF773aDjb8EXup/tDAYS/JowxJdJ3Ij7PlDO
8fdKsONbB5XwGR7W9SGOI6p/GNHFAiVdMFA0GRi4hsbxKqziNnRo/T7R/u53XYAW
QKci9yBffNDQnF/zliG+ulK5kaQ0uqtDW3NfYICKiB/fw2Z0FaM8TxzLEpOEL2j7
wChJvjZqYy9Ls41u6P3Ewf93Fn6f7IT2no8evc6JikPb3Sd2Ka2pTxBRg2LbRgSY
1OdRzwiJpRFu0kIrEuOfVpi/IlLN4L1s9NMeddTf+EcGz2ukGZ/eNbKbOOmSKYup
uxMGXjE1EEbI98JWeiSdwnr8O38tBIueD4/3dFNW+IQKsCaoI0D5ZGRNSUkpjECp
W0v0ErGQ1LsnVe166NNbUbquqfCAZ7AGSTfsXWFVKJhjCy1TQxrHFYmT1HEgyvnJ
jx8jc88rD2sq8emID6V/pikq3pcJ6lOXGtO4BZiCE242hFf8QgsH8ml7GOp5Yfel
f2SvnFwqMq536f3N72MIRkY2MA91EtZYKhv27rjzjVcMG/RCztAWNQnprEOYJu2U
5wmNuUXFDzPK+Mpi0zp8qk+3iNRJIRwKXi4xIDEjwMR1rdl/XyU20+snxGWmI18Q
0ALWop99yUNf1Gdsje3uY2lU8Vvt6s8d/dXGa5eim17ABfmIHaBr9hjJA22CnyjC
K2du5eK5LEMKxz5y5bpbojMltXRmBGXbbxwONVxD9+R71TBZ8MjIhbMfRFm53oRc
au2KZstJfcbLVEGj3kGAPsRkH5nBm5+BkV78Q3UFW3fFKa0kMy4eupy1hTkhtkiH
NRlo30vZ2Xm4Nt0nvFeIFcBfuQqVY5awrUYOBOD7rRm4ixVhfyE1qQ75WUoWUBXp
otb+ET8QgTdDGadO6b5L0b57FNlY4FXwRhI+vvOaAlks6X05/M66nkceFV9jiiFP
q3rCeuTU1P+X25ENs34tvdxkL41uHRH32VZM9UPvpT6RXF/QsrWoMRGOqOn68rmq
isZNrryAMp/0hHT1goqCTp7PvLCO+MOK0RkIiuWv3vjcdZtOEAYmOAKZhPRHp/lJ
LMD/2Qwfh0jKTUQHbKnTUfTb/5/jBIT6ShEROHbfQ6EdA1/QbQn9QKdsT7G3GpGt
cJ+3T+bIr0Rd03NmjyYfBDx9kc84FEiLBGv25AV8y99DGXK64r3b5eHIFUe9Qxdz
z4gp24xgQhDuF4XByJ4bk0too2JhZ8iV3G0k1qiOdw/3n+HmqsvNeIkupU0B/FPt
2CvK69aOMN6JTELdY0JEMNckbqu9DzbMVXWOlw/fXaAU1nILGnpnGv6inDR+cwfK
ndRi/2j87vbg9t7lai48jaAGck0FqzwLheTGBwoJVj7ZIVSFeRabxvcwQz52UgF3
vwkG+E+4km3JMfPKfAj0ZveFdmoI9BpLdpmv7m+DPlMe4HiKjAqifR2jTFol4e42
iC/U2qVCYeaZifygEE5ZGEHznqiCQcOs8w63TG7ngVbj+bwFW9VQbSNwL9s0K3Pd
bbWblwC4lsMiLkBpdtqLXFOTzl16ER7rNMxnQYCCf03ZKy8kNtjaFHoboKBcDurq
A89ywkwVkHnRJ0gbCVp3RiA6Wc8+9awaQ41qwMiN3VqiHvyDMkSmbQHAYU8Zjhk+
Ztacdbqju+u6wFIWa3Arpq8yQ3HI4vYnqJolldstgob+gVJTUIHVBlnunAY7KhC+
KWF9w1lhujkuAgexC71f/q5sqVbDH/miPrLAIgoupaPknTRvTJTENv1q2Owu5GU3
XbgBgSzWXZNR6bbAFVv+hMN+zULMKpofxPKtz5FLyiLAgOJTF3NoGz45SvA7jMLk
pM2CWt0EXuOfrPwZYOe9JfsQr9qaTrHlmuV6IZ0KzqBONFVGtvIMoDOr1udnXUeW
xAd6Yr3ewm8Jj0W712x+WeO/vW4Oia0gU8ZpJOpmm/3bUEks5Q2ijqeCb/uHUzuP
9nIjnclfkwvDSfkeLu8Js3IV20YZRYyun+bjxhunJzIni/xqrnfIhqHLwSPUlc5Q
gsJU83kdSuE2FMY3rLnmK5U+V7MPmCYrm/zdi80Ew8zRV5n0u1R+46QcJ+cjo8Df
W9BM8hlOaTzw4ZpL00lVraUNtnrchFVXFliwg3E7IRITDnkNyz1UTOugirNUdS+b
KBJNTZVTgLwMFSYj5OV4FaE5xYPpRMRwx6TVLAVwLz787/tMoeE0LgsD5Psqxhqz
WAE/ChBYfO+EuiYpZxrX/G7gOjJ/bvoNGWQL25CkHYg8QmEA8sohSoERUB7Mqoyk
2lXBQhah4UdiotUKjuRvql/nl1H7wSpdQ7WRvD5GjOiP+DGewpR9FrE1JhnR/PAJ
JdTOl7G0rzCWB9Uli27lxWCIyXgQofmUEEUQd0xH+Po4BlEn5oCPzlDoJPPMyX+b
Vpq/bILP2y3EgNX0Y1vyARiqSNpvXfi7DqYWYLTkq0HVZt8sjIyVF7NeE1ZT7HmP
9Bou02O6t+Qfc2KE8FZcSRb4eHkZTsYOS9/rwudI8fN0ZAfl4dRFi99Djzq8lkLV
giIC3xpWPOLYJukOYT/eXucbc8Jmc1NotdEPbuTu/0x31XUmMFSmlObDCYEnwdh3
2BpPhT2jegFyiNC/QiwAvKLwM++/0mK/ye8OAc4SX2CSgQikiEZIsA4k9zw7kFk0
lqwwAISmXx383xBhLimA6S+IA7r2s1iUom2b38QhVLb/SUvLl7dsvK8hjaFtaiJu
ALXC3/qp9LRyJqeu6R4aRuVrrxnD7z0ULlnusIvHW3F4QsC6tuWWidO6LJTkP1K1
uzdap6JR5DZUZtKBejcpkxf6fIZJQbfC4t06mgQPPBNaiXQe6ZbsFY2PaaKuGab+
Z/APiPxMV6QOLm155slgQApLQozFOGcdn+QL5HljeQ9d84LSBO3SGxdJASBwQurG
4YF9usdMMjFv7EfGDwzAfzfZ31oTrePBJv0SEXBoRCF6daQo6OJ6UZrUOJDJv0RY
Qcjb3QvIfZ2c5d5tv+ytwQzd4/Rz/CPMfaEBp3CpgwVDLXvjxMkk6i59F5QLynf6
xY4122/RclmT6pwesregUXEWBYSJAHDqFQViXHIq6f/uUayYFJIHWfqgJ5zCS6Dg
bTnT1aA1ZpzG/Fj9zKL278p7uOiM0GtUeU22qI/Q9Eqsl0xNuXD9JAYy+u4Xju/f
OgvUATDaAtmzgrmTNZgp6DEKSKyWDQ3D2COagNSdDZWV3llOYdMK9G81o8JbtGfs
f48KKQVxOijXUvJ1zEqPRHm5YWHe6FkP0G9KMlb2R2IYQ9M2BjvqQMhzo5WwWhTz
j7/v+I8VbTDK/TUKQMtxCXxy8lQi33OEnO+ANU/ZIjv0szgbrKzhvKN6U3eRdS0I
RJ1TxEJYmKgDf7YmHLnU4z7HzVuubRC9Gc9aaj4KDP8DRBhWK4bH39xjrIRt+sOd
I1DxFTzaWERXMV49r0EAjWkxlPSOSTUOFAdrnPuTcmq7qU050vEeRHbIKsK31Sko
rzvLJKhNznG7FvWWDP5+tsvSP5qtfCClCqm4q5wISMNOYqOwjIVD7c+R9zvb5ig0
hCxRhcwBhvIJnv+dUXi2BQhw8fa7LIfV85tLpkwXb6ICdX+Xn0rCs6jIGBETiwjR
Tlq66XC9GP9rzCgS8vtUmFvOkr8i1Vu2ae9kFR6U2VYMXhXhQzRPM5lJGc6M9SfP
UMA3UwHldrBgxQiuDpJTg+C53oV7/sUAID5ocXoWt+KXeoQYqMFVglDauy2IpNRm
plZZv/+ZuEJ1YWAmm1lIW0DokiTHp4A3NA+Wh3YYiFIwHL12jnepFaEyXSQIrJCK
ZrGbhDOu0nKO9ZE7zIWnOTxoodUHvFLPz54QTib2Q8C6SMHbfhbJfptoZ3paleGo
XN9weQdlef8pK5K0GwBoKBAqxJf+LLfqwdhL1FuRsjSpIgERnC95sAlr+F/qeUKE
xsxIPDtiH9t5j7zSC985npVjAfLpvsZ6+P+KlKhTiixVyUC33qnfBH1uWU/iq5BH
ARVZvqLbG0s04r5xY6RvlthAVMBG6wjn/FkfkMJZF7lMvMStRYwGQYOACkG8sfwo
rrcq/SHdN4guykJcvHnLSby/vFs4Ey4MBWVxGDB0mbxVAwRnUURcjnlIlyeNPBlA
5cpIZXQaVg2d85c+YTzINb2lQVA9achLAqPPYTqRqyXLwceayQL5wl5nsClczF1G
Fztyu+yX9BrlavpDGJx2+uWqtJUUQ4d6k2tj/cbI9YUa1CuDuBvhsb/VHRel6Gya
wr4oU8UQvG2xm8YlqZjNSqjSnL8VrtMdMNLJWP03+BiWU2Hm9e1KjWHU49QbttYc
+mm/bzLgBpQAp2HLJw+MA9ODCH0wO70K5JvT2dECD23Z+ULZCqB2uHYh/VpsqJ4t
qTW/h8RHtGewCKZ4L479ufGjVIhYjuGx1EPRNcdc65Md3l7gKEqlLjsGKvnBHw4B
A/MUDXkAgealkQTWyGGeSEyhm0aeANuYd5wt6n0Jv7MqMd2xV4LHbQPcj3IIVGdV
ee4Eb0+6MqGOwodlS8FJd2DtlU+THsh4WyUryc4Mhp6CZYCm6kMhlys1ZrN4WOnH
sXIYX9MAMMrBc3ywRMO0UcTCs1vaSEAlpxAThtQlJ/c1B3YZYa7Hg0D9e6zdyVLE
rwuBtA7D9MTKYRa2kq6XGYE4+D6zbph/9BvCOS5V9XvLWvPcKX0Ll1aLNMZqbvkD
t3QUN4C4/jpQysenSKKYm561fAs4YOo0Xbgb1YjsIVoPIzDJ1uT27qmvXsMplQGt
9F6MgXujbKtgw1Mc+qFx6PQdYX6DnHHvnP+hKq9QkC0LVfzlS5V69M8DA7K1H5VB
d5PRrtQmpCABEMvEQlZokipPiHChEZ5KVD0szStLHjezayEmzwtPpUPDdL0WcfCx
Sr6lQvCYqeIe1ymeK3SofC3LRTNhHfXxwzYyFFPFGTQClr2CL7vxk8S/JbZ9mPMN
J4kYNnwgetwMAAQZTSzHR8o0Yg9eK0fXAKFJZEmb1L0zy9fZuGsNv4SiMzXejlM/
V5HkDKCT5Z5a+m36Fhmg7wCZJ7B8DPE/UBAyxUQCHzCahbehaRejkkUohOlzTdhb
8XhXgfKAKeFMCttDuUPk3At790RIDXyaLkt86imP1DpBNQ7S0wZW6kTmTYVg6tMs
Sm3rOWVXbrx15P+qb0yCI94+FHGd7m+irvek2oirWz5yC7m5AQFD2ME6kwq8ZHTi
fj/LC8893YpWVUMNtzn8eWYVpvbOINDLbWGlyqoUOxXWpc1SYxck1sZ8gR/OfqVW
VyisE89Id9bRkQwzcmqzScW8cs7VzgbO1Y3FqMOEmkjaFvEWWT8+yEZPy3FFELFa
3bVDkTSDwZ7y072rvTJ5LbOpGZg1wCW0Sy+os/L5LgW2xO+uhCMFktBtHt2pPvgR
7Pqs2RbNKdRPWGhK6+pfO+NsLnCwtc08DC1BK7n8Df/flyTvV+MMeLCixya7nc17
3qbycE0LIhBmqU5qwI+PovjOR6bnR3dOk4v8NV3R8Fk2xVLMlePOVrEWzB2cl1qe
8+y/ClF7zxoexX3VYLIoycm+SxViqyWym4plHLJHDq94f/GL5zojuQgETQqY5cG8
jg6CoXSpTgbsWyoUKltBuonX0/vP3Z+uBv9nj7Mx7Li+5jAinn4Kp+BRnWa9CWWa
9LkjtaGz9LDvXAmgYWLOSV9tfSfkqmUd7kF4qZOQvpQJ5YFAR4l5MnB4iVNtJiPd
oSZSP1b8pRmWy0zsA8NmmsqB2OJFW/DdQqCiG9QTRa9/SZ/Ps9ds06VfG5rZBRBH
Gax2IGSG9vCkM3Wcv1KlgIqTinAxgQj1+lYFvGJvgRAUo8xsaikAoNet9fhB+dTV
LUW5mUKCEWrIxpuMfgSRSvN3ZO6SGI0QjbdcqnIxxbsEEcRRXZhH14ap7E2jWwtX
Nzug3dKLYr9L+hKhTJo5IDrFetf6mL53joLwVHZ1u7YGIp8cOA9B6Hg0CONPWeo3
COkS9mvi4mkNWRSwkeiyHVMf10L7Yw3vm80amyhAWrAI2qIGjFlzHsPc+/aW+F2K
AqqUFr9hGrrRQQr7AgJa05gOaWAHm4NkI8Aw00QXArElftgSAZrLYVhAa/R9RRqP
/5rHwJq3KeNKj2VdMRfYc+FjSJpN4adScA4LZwlyMLBQLXdN91ju1zU2KFtuF9gO
xIMjU5829IZc8GORgqLwNxiyB1m6Q9OWZ7X8tiD/cte8X3IaX6n31lFGMo4AiZHV
2idkD/PCe1nz6tP6w1avXWIM+zHP0jgPvt7TtApiHitx3F4Rh9aoMBLNMTDPCBBI
IaR3Ue/hS7Lekdc5cxgR2HuEmSzY79w4kcJH58hHJzyW0ys8hXS49YQZAo4LpUgO
1ie2uUt34b3Bkvt9zox1UQuj83oOMLex2u77cwuwAx9JL3j1mXLMqhLOaE+DBwXg
ppoOp00bXvAkIwyCKlG1q08Eeg2LH0c7tOZctTUC2gUkX+fMjW752MZxeSo+vmwx
7d7oxNiQDE6q9wnO570fYjrt5LE3qmFW8ExzfkS2Xy2wcIbKbR4foTCxuBbOHe0x
luwi87LR2CD2B83wAVhMxM/nNAxzxjUBqTSOmfG/h8G9I9vnX13MzxoNSFQD76MN
90L946+E1EavoTolEqxUkuEMIli+oFz8YWEIRumLG8UjYuDR6v7ceGyuiYmxyRTH
DUCX1oMvAmtYp7+OSpT5eIwP6Vx+pfqmS5e6I9zQYHBDh3JoXkQmKEHTzQSLSWX2
XH7nS0I1msJFtbjD5gVWBK+RIlb52z3aolUNrhOZxoXpz+DdpRFZEp53JmvVdHxT
ljKdYxatywDBbSHfrnWnNsPiGnjivooSIBUco39CsM6waBF2Rx89tNpR3esaL7kC
pE8ZuBDZPlaCQcn9hYsPcslpVQ8jE3vvybbI3LjFzPZ1oMIDZSK5T2UuLnKLsCcM
ROi/rDCSJo1pn1L1jD+UOgDVV2+w+Yz9Ev+H12ajIDz+SmjP9x28Fj57d/nxOTny
SDFYMoJc6r7G93jAFT/k2Y1WK8h+tNhZeSXEx2IsugK2za0VFSKsrbW5xa99fvhv
p7rb+XJaMvNtvUPOCYu07H30LViFQtcYi2B6zlUpGkULlUWbjJ+lwzSP08ah07ex
1rB/8eO5siCiZ0lPwP4xjIOlBbBJ77+QYG3zb6IHEEs3Nx2YhIviKDXnwQcH4eC9
EZCzgC4EQt+xLfEpw3tXD5RXOPssX19aVaFTpQNHzAiQ+3xEQRYt+k21ErZcrp6c
6J2iWXvfXj95oyuRZLdDBS7s/lOxGVOTqXv9E7ISjZnnWO64fjta6kG2oijx7N4Y
pCpAXkdbzE1qhjSq67zrkcScpiMGJg03SChHzUzpYGu8TnqbtIuUvbrXCT4cPgcB
y1uKwpWy2Y5m3z699xDiDMAt1qMaca+Tl19iTe4rnKtVfDXjdb9B0KlTl7KK2EF6
PsvTtYdFpGLSqdc32Hpt2bXUyKFfvOHck1sKzWF0cttVzTnlZkIQG6cWRqR94G8+
OwZYgySwZw36SJX+lJRdftbnNxj+8ywSjlOx09cv0JASlb01Qdwr49TUqNO+Qn4e
DgSDXKjmMuf2NeaeCNe3T/vOKJwvrD/y2ns2PYseaPK+Yj3fSPPE7jYm9P/VVEwH
vNonBEqjHKC0Dr8YRqVmHGbjF4WNOLaUrAn4ZBmnUVTMtO9TDnWVmSO6+gAAVn6e
iIVX0Vs4EaZ4WgQktchHZ/u8/MbNtbn7hv7E83Z+qSkIgR9zum82XlqKJHurpcd6
olO+nazuNFikJBcIv6G2rZhzE55nliqvXvwpe/QXWDETP2sLK17/eeYqKgmBddIU
xYGC5CDVnIJOULTY/E3M1BZsJa9Bfh15lV4FJht4q5J3/DBCXOkCHvfP3Gdtm+p5
X2rI8Dd9Mxp9ffdbaWYhEwdCuJGiO3zHfVI4vs9Hw06EeLaPDl1wbMDIYzAGuFsT
FwwsM2DZR+dTa4oTz/MtHJRtuCiBsPNZ6TAriqrQKBq4wPSZAux/j6HuI7rT+/CC
+qJwW+cFfrrXU2Gd3Ss3maUKuvKmXN0znK/+iIxqwwWbsoR/EWD4fLoe0to7liDj
0kKZX2RifTjd/VAb/pFPwple05+Kysi8eFrtRYt6HnXQc607JHlFh13XsOe1xnC/
3it64GYtEAD9VOxS0T+owCt4tTHf7Ki+VgE4khaREESr7ASUK8AZAlGK4gb08OsQ
2GDm7RFzwjXNvSVRPm98TSLmrFrEn3LiNEVDtV0t2iFg938JxLrh5zxQE43iUhtK
FK9sBoWlEIFGudZyoQh30rrIK3T0rhQKBxQA6N0jjMpVgC/kHJPqSbps2G2Dlco7
fhy7W+LeY7UUiWu1Y3imB7j1nz4B90koJ+IgoqNyBXUulbL8so47FwwzrvqOC5RA
49tD9gbCMDVRfi+Svklx7LR8LF2c8Kbgx1sIt/sR/uJqPF9vUQpjvV+HH7quV9V0
YB4m9azYQMzuMcs1IKGroj1RG74CRRLuxoRLkig5G9IHaVnR2Ugz5OebljguXADv
rCsaVi8AekV8XKyvc7Apg9zwzjUh29JW2VXp2b5uV5ogaBmVVmU83zsT0juNYv1A
IGe/nF++NHxKzOUYmLpf1cnZRzUbYVUyQXJ6T4ZJGvt3Ayt8NUW45hR50gDNpNxV
2Q6qgxJm+qhJy0RxSDfTEHjndvceLFFSwP6xDtRsaDqg9jRl6mmKGeDKbKPUYUjU
8AJtdgQ1dWhdt++plg4p0pp88njiPKPO1cMlYWE25QTfL/JzIBEEiJ3HMR1RNpnH
WBcTMWVRMyy9/w/4ofaDSekERATspsIv9Qq3da//TY4=
`pragma protect end_protected
