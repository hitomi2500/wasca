// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:33 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UpVruHOuDJzGwb1gUw5/NqcuTcciJYYipCYMKsSDv3myoXPgkiCtoBIWc0PPKIOu
+1h0KE3zU0AXrW0Q8fm4tcDYB+kvkEeStb+b0BLIjPYZUBcu2QXBJnlRmacnb/et
100sEGocAzdpfWCb7aQv88Qh9psPDdhnDTXpc3xCO4E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
Pf7Yi6vd9ovQgYzR4L/jCsAPExMFSSWiCZE2AKRRs8Dxb/TiIUsvuNV3OcKZ24Bd
QvJ2n+OG6/mKCutuWahPhNK9pQyrSqi5cjrs0orc4qkdan/5+Kvf53nkXfsRxZqN
XLMDZZe+R06uZPg4CCAiVrj72wETVFIo8K4D52kmbOd6Y069V7s/Xxom8pojZwXT
UINTQZHEGEjML+uYAqhHyQ8cYm9NEzH5ZMWdbJdyqZlVMAAx2rXS3RXzxsrJ4Nkq
+KAMzdUG+uw+VGiJQa6r1zKShMVAOOV7pl9csRTCCyPzkf4V/dbOK+GWb45cC8e3
85r4/+2ME8MTBDaGHO8jyAxcv8oarUm/Gf2XOCIhBxbaTjybks6FHzVTVOeIs+kw
kLQrXvDdO9Wj6z1R67rm/kqHP4SvNem7Z+49YFM72b4R/SThNbYin9Mhp36H2Ilj
F+Kcmm6CldP9TwQ2t6VLQ7RBCJweG5Tr6h5cjvonoSwpi8dBC1XL4UfofyjhZ1EB
YNyyPVKV+ge6HQhpXZIXzShZBAhgfYK/KfWysbuYyDBI2vpiIafjezE0jhZeFMmI
amq1qYRBn1N5YxgQKVydGr+ucvD4WCkYD9T5q5gxdmRd1haSUvYjhbXPZxbyzJsg
kErTG5ZkC/8wKTGuzIdaI8o/vHmTCNnKyC6aLidINKKHocLNm5aeL8M/Eee/nXFi
2HLNi80dfVp5JVzUgjjr08He65fCHCGcYlx404M6Go7W0fKCLMLo1KWdoJyrkJh+
iw2XE7vZJ34FQymHizWy7B2gZRUMkVSLeIJLl4FLELHZjBsEE2dPImiHQZDx5//C
y7iY5DdfyRFIA14mvk2DwG4n0KRiqtM7Zd1s4CXmV5qofkg1DbGSx+uRpL4jbzlM
veQQfo6jxdVwwtb/OskUKEj7wUT5/jYBVH6RG4c2w0HEQlsevYOh0JYtaFYy7syt
HeLG9FlnAiod9DzZqXqbv+pusIoikv+DdjFE6Z+cOFQahazHnXCQsoKjMwNMGD8u
OZitmXy+FsOg7ecDxIqbE9PZyPHocU2kdEN7P1wERXmupO3Qr9poq4nadvVWBaMu
7qSUDiUux9fcS+Q1AV6jz2oNGq0yqUYrAlcK/dKFj4+5MyGkrThE03QY6PN78HRB
igmT3qJq7Jz1RmpAZl3YkHH8qjlo0zXW5FjzRPcV7xb1IwtfABK8+b+22S3pstbE
BObf1Xm8SDg+R8UIBRr5ADjLtSZLZcHaqAnAjwqw426aDBF0NR0u0VGmJ0xl7IfK
DmdMvC0XyvQMRjpEYnTqv7Wmyl5FfasquXLpV2gS/GvXazEAP+sjguXJlZ9LXl6C
HeBch9cFH0UAcut2LnHJy/rsXCdIb6zHabuF3rRJEBSlfwnQVJxGI3gftEMnNyUy
udYH8njQe4irszu7IzFiVADYTJjskn6S2r8ywWs29ZiOb5EH8+FSN2UMGkXXe7o5
UsKIYgsUO3m1NLtmRDYH5jpklMy/hnFzn5lEDcHk72ldem6TNhnNI/YH0UJwiBG+
IH2DiwzqY+LLFh9VMe5bg/1Jsd8regOQLg0CeoZRgew/VF40nBTAIDNnspOWFuDj
Gn5CzHhaqwpl8OZQkxzC8hN6JpLeiqcG6WyudZX/tTmBpsp6a1h5FqwYq9oo3pIN
FvRHlFyDWtpLdOqFNtNQyQLf/SKAT7WjsYT7hMSdncfDBxhO82nYI00MKaEk7Apu
1r5J/Zgt3L+pstaLhE1T/RgSD6ipvC6Ek1NKhLpx6Wps1Ohc70yqdCErgRrfyWt4
hWbKPRNyfIiRl3BP8FxVubJK1vLl5F2YRfYTnxIvTgKzA8vuYT5sr8UTDY4H44Dp
HxIdh0Wu6hjHeQ+tZruqLY3zo4o3w3rCbv/HkdjTg7UfiiMrGIyI++LylJtYsYxM
PcrdNYq6dqkmknrV7zr+RUYmKM1Hgmx44O4L5Gj/d9Ai9p0zLpgPTefgesPMgnMX
FtCfOPBAM2G7T/kMYjA/d6KObuWD89hioaJqFa9TFczvCLOyy/8qh5hRYIPyK7Hy
bd7KBydn3V7jNNaao/SUq1ZZMRFr/tTFAvl+KDq+VASn7GnufVFJAxfG3GNw8Fb0
o2huOrVUw8WTwOOFgeOISpvGLtJ0d9jF3h/iSDreB+E83ZDm3QKQQS0hUs3ciBh1
EfXmf8v37ALeR64hYdT/OHCuyL/Q08haVH/npmPm+nrYjZ08O5rgX1oXua8PuDfO
XDSjBTN9mshPgFmNcPysvVVKAc7UNKryFtLu3QXPt5DOkY06brJ6kvh7IzxET89Z
pi9pGyS4x4OTRzfjh3yMN75tCULW4csiXmIr6qUBedB4qak/Yqq3bvGa9OrRowXs
eS+dCPhaDuRAQhzuhawHdlwENDbt5ClkT/SnSOHcIv2+VbMED0y+afp2KMHmQdx8
rv4vlyUPxeGArVwQIpx2LzTqob2iCzmJEodV8xAADjrZQsHoyGj3qyWMc72FpXKv
g8HwJPRDZDH03vmUi/yZmqpI40A8pQdZCxualJP8IelUfv2JzL17khOY5S7RTmwZ
4X4+1tJgMFWS1lm4pbnGcxfSwQqSFblR5HYrXJbDDsg4QhGnC7d07SMDdv9ei7jz
ZG14kKRCnYjKz9kuk5V2jhiPYdiswtydckF5oJQQrjfoW25ubjqm4yU5fCh/MYEr
j3OwIkEColSM1FclBnLDbIYw1DCd1r9CtBd+zkF8EqJgkfJ52+yhAppXwc/RfQX0
3S3a90wp95BHqjQ+o1e5QAKflSi5AmOkoQGkukglycShtZ8MgA7NeGxmKLwXEtqF
jdJSdx/N0V53eiLfGkiHnRXx2ZHzVZWPvOa465IiKkFhWM4jJiJj9lL4UWOmb1c1
VcnbAdAlUOD2lFI4vW6ntKvKZFFWCx3NRrpWOtZHoK2qKHtse+TpwdGJjp93r0eX
JWlxOUGpGQ49yXdYJtyPR9Ey0X8SqRp7rhFOXj1LBQMVOm6ByvtB/o4jcEji4szH
u2U/vNqaHUCMGZ2i4e0EnvHr9wiaX2yO8SMpuGpP3lYiCyMhThOpzobvUt4s8Ca/
p0bJaGTH7YLGvfLEM1QdkqFAi/E6t8zEDW+HrwpQDFnA4WUBdY1rItMbUQe7K+gF
kc+3aP7rTK+VAr/VuXtei75jV6J/NJR6SBNtMjsMG+VFbf7wUOsN+nRuFgVOxEyq
a/2Vc+p8efwDEIpGs5K866IdMPACr344bsA6dSgHxoC4ScLVyqLocMNDJP938tFT
qGTdO9KZvtx/NmPXEiBWXMiUY1BfIRr4nwc8ao7uNlQ/zvBx6zONynVqNusA276y
+vG41+NQIkubWjTVMP09NCTMu9x+XniwiCaTicXKpRjdbbwSEXECDbPu08XAn+No
+XoATLwlrVjtuo9XOJ2l9O9isNNkHy1xiCVci8qmkcC5X6xVRxTN+A8weKxcpW5M
kTpsg24DjBFJmJ6vm0lzIsXqvEV8c7TuBT//9wGTsksuQ838kjjyj7fwXeLyrl+t
OrNs8gRLvdOxPJPoW4oXwzNCcJL7X4OxMdvC2RfB/EmyeRWBpdNjw6w/mLAIJn9r
yDLHex5OA6BDvTmXIO9UYr78yPAV8MUs8NGjD3oRCFiulD9UajrQtbONtsMXv90r
Q74DdZfdUBg3kf7zxC76eBwRK3kaV6nugEk60FUNcsxnaqts8NaTfa0ptrqk/15I
YBqb27OimTWWNKERCy+QLV7u8ETVTgu5x6NnA3Q9xTw30o4liy+yj6BD1X8KL2+/
ikzgC9GsnMoUivqOTUrHXIY9vZVzR6sYSd6lxyazkHo7TJKpZxCNdv/PAj7YWni0
2+s1eq/sgX9QZ3X9Zvo4EcHBTef0d5rC1ddSLHbTLCO+PEqX2eMPsrKfC4JODOsR
PpMpJPe2vq/g7lYM0rFlAOYwaIe5S90iofgxe7f0ClQYncyE77BHlupIrz+XszY4
tMmlXhbgRKAJASoDJINUlx1I+xn+v8juD1GPtkVk+cfpgojSgC7N4FuBYNxjUU6I
y2RHpWmtHjlsL90Pw9yCU9ySORWOeBMkryGESycZOfhKFnT55CLX36QAyg+6Oags
gKWVc8thROh6VNF5OMGWr8bKumhESxKU2K4ykmqWEtp56gPmJPbaNICT0ufQD2tF
uiK/ujGZxqxd7cAnIYNX8Kfy7jN4Wm5q3dewbVZRGX/2SpFSjz6F76gbm4m9goTr
FM6j5Ihi7IGu+mQi6UKsfSXPYYbWxbM+crPA0WVZyZh1tGl6NT3+aVOAe5i92fMF
D7VssSSxZETzKZqgZP20yRNcfn6XZjbDIRUbqsIAqmRHB7knwVhRYr531zMg4IRQ
JfXGdN0LyDrfhJkfBtkMWeQGU8h7/SfbOWn4wmhQLyzbenKdl+Kf/KkKRppkuzZa
NBsXT8Fs2wQ5qEhGepX/Bcm3CIakrb1FxnkiKrjSPaEA9yYZO0/E2R0qU2NcHovE
oMInboDc+yWYyAVWIzeaAKwRpxYsFme/snrG1VOliBqrqBFhp0xs1FEQzY7r6UHD
TKFbl57aBbRg5Wd22fKanySwp3llBHyPouxBZqIgDlMYCC6H/C+4NeekZl0sp2iX
7g9NBlXQYsy/UWGeLbmV6fz0mHJdZH1v5y2IDA4coqCjeTdB2IDt9wv/FVfp4eir
hvYam76Sdjm66sOla8draMuaYUGjzcRVZlyJINaHLgIt6vn3jW5DIF6ICvEU+Dbe
UKuCiAMFIkSqIjuZdDm+seCCBp+vQt88q3IvsCxeDIoXsE3V9Ee+Cxlo2bJpytRU
6ZPHro17zAOO9I1j93osQa2D6qgmUOXQKxcWyRe+hOwuE7B8LVmHKIicDhVpodxm
AXzMv16f3TRfbTwtQe95WlsLf/SA375woZr21UHj21JzgkjDbMPDE5rUyRf33zuz
Jxiu4qwB2NJQGOTwqZ6WksCNHu51VkOwgm8XICB++7jKl/j65QX3Hk4yWmEt+wYO
BsSzIotx4HaMoEsgdFte/SdL5WERFX9zikHa45gy4xY8GXZ64JYuTlamJpM2OYIN
Isure4RWApW/4sW5yrkbHbmzU8UWqxw7sAToWAs+Kijg76/vUTf1+vtmJBttf88V
OwlDVuGYVhJvEeSIHXJiO7Rfyl7wLXHgQNt+V487gqqz91+fpePbV6bBMJFT++N0
WZWcJzTPDs68MxeVqsn3D6bbicZ9ydmRrHQX9WapZ2Hf6PDiYxEqQWWp3UhGTSAv
IUuCND3fHG4QRUBis7TTCwKdTEt9hULj1steoApZ848JzJ+fl+XiL1gS8+EH9ozf
e2zndzURLzWdQZamXziCW6Sn4lgZT8fyAJSHn6y750NXn3M3v6M9aeoGdI6TzoOK
vCo5SItXvnkIZixpxBgQ8ukrvtdCnkEFTCcWH0jFaaAQ4J9GLEg3VQ62allY2s6U
XSLZGau/Z2j9Te0KB1/+Sz/deOEtbgdRG5ZSNDUYBhLdhY+XZ86BHq+G0Eyf/Bgw
gQbUCHMhWjd0LLnpcUxseXFFRlZpNAxF/+j2D4YSqE4Il7XR4YeBLp7jdRVRaFkQ
PUqV9MTwJr+Z6iKsgk2t85RmaquqnM41gclXn7MU6EDXL/QYSuwYV6QxGlrP0L2R
9nkxcd8Gw4YYw+sOz58EhUyj2b20oGWwd2rUcaeql42wLXGL8t6gZVMGX81xTGFj
QYnf4PyVrQbsz0SjnsUxzMk/C5xWd/fkGue7Md5PgS7ycAWMMeyseOWqgiVt1qnE
jdceukB13JJE+Vvcej9OAhvHxpxO7ZDJLW2atVf0FmG3J51Qmd8KUpZTgEPjdxbS
xkgNFW5OLDL27lhgwpg9ghwIWaiW0nULBxtlXn7U36C3Yf3P93NtDLTS4LX1YsVT
vaSqBuQ0KSjRSPmR4j8b1Tz06ws3QbSfa0AbaAkQFKhhqCQJ8nYTsUzY3PGHt1ac
puoMaiLy5RssgQJ9zTB3ErN0jrP9+iBhR45RxUtyW1jTrxHTJcBEyPFPcq3gjVFc
k2IT/7+YrtaVleEG/xBgDssMWuhQo6TGWw06X6E9BPfxFQiTpzzY1+MaOqTMFN9z
DrVjEIxLCrs5zhCYM5dPBBGwGayenX+af3UDuMsaAoIs/b1FcoWBOxBC8RnoEyv8
7DTgc2lS44nuX5gJqJ/zS6F9JS3XNiQtwAF9oykcw85+v26nhMBUrfdRo45G2LeB
edqneHbrchI3wVRBPzYRRi9NlZNBvmRnu5olo4SyJ0TFkj+UZ61pBSF7uOvQM9e/
3noCchYMAbE+8YM2qvJgsA/gAgr049RDwQeSLJY5EfWvwwT+lp8gpImO8U4usdj/
NWYXnjEBAAvD9+mfGXwOKC4e3EZhH9zZz6VYaHasYrgobCthW5r1aZsjAWCwa+Lx
AP+CdHORvyte4z/T4HJ0ZKZbAunTbDb4FkvYpsfCEetloPUP17f34cGhBEJ6pegj
G+cQXb6V0BPkUVCzh8zzmUVZaud4xN0/LbNbr/3ExTw/F/8f/dnYptwZ96yjX+ro
ettdkxhCvPzvtN7TgF0ovjanFRcjLokAVxpX2uVhJMPc8DMUeRYKbP2ow9H3zMuf
UPkvsgkNs3/fDE8IUGmfVA2O8IdAbyMQjw125gNjF8Luu7t5ZsJG7YqOr9V7DbOY
wZaa9ob4+kY7ELfVXJlmDWp7/AaGRbu9gWXW6vw79haH+rQLGZHtzEHAJ/xScO8U
vu5Zt5eBzcTB9xshKTtNrBEeP/cseb+BeFu8owTIDv6zuJvcdISfsO6aisIKiC5i
BP/RAYcABgalMN3iuyX49pPV/ZLxDuMKVKVGDBwXXtUteSPwwhXIhMjBYMtOdLpd
l2dS3Fu7DJBFAFiKw275BSX8EzQZgrZhejnjI17GdcdcaiPN3PZcP0fXeRVxjp4x
ZR8bY9RBJRfmZktnjr5tPBhEGy3yNm4bBhrQxJJGwSfnJuYK4RGr6gPbcjG4xHoY
5mW0Q3BlzpU2WKYELZh2jw5S9/Qs2svQyXE3hfhyOHA8iAFpMcX54ps6sCdtsIlI
6esSmB9ijgfj2B02NDq+VYZ3zvOeFVDTqkGJ8mutbMfj9/OS3Urz4XpF3O9mGCwm
r64/nB2H0yIGDDI6lzFb40ILbbRNlgY+zoPbmIBjcWjJz8Uck7yjk5XnfCGUBoNu
qHML8G4Dl/FbaL2nFRRLwI0qCmLLhm7NaSGuo2CrpfC48C+cbAS5yV7MPdG/xRoH
Fqta7soOfAKISFMyR6uz+LmXONbp+87HQp7yWIDDc8ufN4LPhlyM4WWuzkwZxnO4
hOG42O6sOZGqaAis8PAxqyxBwziaAOQLJE94tNhLsbwMpW1NbCbrN/N8hyhXdjHN
nu3mlhavDs5IZd3xaZZ+6I5wL3uHZg1eoaczROlpJn0rmb6KjAsMNr8ZoSAtKJ5r
`pragma protect end_protected
