// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gZxOwEdNUpGmJInzY/9XgwOtVQtDC519GlsJLDvqn7wWQOuXhm2dNaSytk4pM3xZ
FHGnanhUH4e1rjxx1bpJ8jMYqsLEsJfLyo9KsGgfRMEbFGjTf9gQ74kHWtMyIGAx
62one+3pkPAYJ0CX/zwGrogfwrcC6wtJjc2WyRlE3bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12256)
5vKdaRqZXmxjH/5fFtK+irTruIXfr5L/a++5FG5lCU/YnGbIjOAmSKh2pM0YqYYe
JkIjcTs8QIVt4T843thiWF8EukeS37Sl3Tu76wCBMYM63ShLztnjobEkj+lYp4d1
yKfxwj9B8Gipz8g+7ccQWxKU3bfD1j+Ke5liapMo8JkjtcYLzwWvlmg6EzTEweR2
iGPMyH1/VtRFow2P41Acbu75KHMa1sL8TqIARlHDGoQHgtYSS50EhLYGm01LhVJd
ubQj73h7DSU4YTF1hdajL4d3WySrXwcYRTC14GuE8nXBydSDnNdMFCO7qsb2vPzO
qcaAK45T+iQBOKOY50g+HObxBKtOHoU3vdcJaaFVv9iOp9BlJo2j6KShko5HapvI
1kIEE9e5HYoUz3hXJUwA4L6QW1RDxCanloaVbjjDCHeTjQwV6HHvDYLeG1dXVkF9
tkDtrfWoeaHgpRRvOtelysTL7XFGWQCyGG6OcIepUIAd7NQyGCG9ytjsS8hG3Om7
5GPJghVMIVhtdsM4ut6/XhSGGeB4kiMjUQHhC1DoHRPUA4Od0P4QJW5SmMloPl2X
gtbHoVP/HTscI/IKMLbgBnkxIUG4DYlWjpMWXvK0B1eZ5cwiEYp5bofkw1lE8Rsw
B+pzLAvI5e8NgnE/RT5hGCSGYwCnKdrCkaUcll05LntS1VxOIZu9j0tW3QF+gsdO
524T79long5cfeHaDCos6xnNX3OfedWQSVCslOqGnIhTEmSt948pjk+1N7jznNxH
icXON8b7Hy6uZjcZ2n+KdSFYWiU7oY6rnegkhnT9eQaP9rOvsIeV7HOs+/U7Flie
0LkJM7osOZnuZEGrzv9bx6Fcqo/HdvOjzQXoU5uc7ieMMnRPHEQWYTeUcmjuYxI4
/+z7bs53uKw2gXf5W9nCOUF73RFBffZmBf1KAfMCjy1Pc81MDs1zk8Me3SmMuC59
j7I75xIlUgR7Fn/WuZKUID8HJfcQJehE7UUMJx/mCPU/xu3zf2cF2Woe6WDthT3G
kE4XcuIYhwPlPvxis37lFFC1zCK1xBW3QhU5sXhLbCuGUgWyjs9DXiRExlex5nOo
LjkjUUva0UTMZIkh9CNVFXTXQLCVrbxrAgPT4bv8GY4p7ES9v4Xre33hyivOtews
kjxWINTVUgr/TKObGE0j7487P0vHtvlTGgity6NY15UdBhk4kAnX14CengSQ9K9R
0KWMNPHEml7iLI49dCf4E9d0yyZyK/uVNJ74SnOvIakBe0vw6bBKvg67E0d4pk97
m46c0JMQI13y5qQfvRg3V2OVbquXIGkjy/MTqElPQOPHykMzierY30PF1Um23kVA
Mt7bLJhXl3n6RbHZBvwZ9KnC3xvXB8sQUAmXmrqifJxqNvs8xDOau40a+tGT2N3U
hyQMHq7QJaeDt6a3amIuDbz9RslYoUryGB9t9g6nNkZrdYYYF+IOsrk1/lZauwCT
mBcJTcgKotFqC7TIlLWvK1C/ONRjZ3OGxn2FSQEjve1E9qjoIu4S+uKMjcdSzPxv
mb1uqZprtXURx9yaMTj6E/44RDwhJmc6d/byVeqo+ECeZvwid8tzhNp1JMQcx0D0
W2n1LyuN3actIutgADy7clfuBhyqwrV4O1VZARnCcoOycVUYOhioxJZ1/d3wFFr8
fvjSjPUpjvECHbx0rf6EiiFUzIARN+ijartYHOALvkthFFNsobUtv526iO9fjfs+
0FhRMk45TcxzKfy5KhilA8NaMzfXDa5tmrWPSreW0B7so3KveRJJMZOSnD7l1Zc4
mYXJJU/woOWE/q2TIRIzXEub/WuGIwgyikG59sFz4N39P0ILpPqqeQ7EOe3Ljpf7
2jTYAWB8Hf/OzybY1iSxybVGEjmIAj7jxVqF97HMBYQTTjmTaynqAFPXcJEWR1TL
DiHbOdkN8rgg27tPbMR3QTL/lTVww1pyirT3jjaFeGrwTr2o8xtHDXX9fz9rKnr8
DPaRkZesisd1Jr/n4uPfJAbcvIT1DRd5ASKvfSa4Nhvth8wrp+xGxWHQxG9KxC/Q
pzVmn/L3yncPR3+kMTmUpPNo74wTr0odV3Nl0Lh08O2IZZToM1JNBsls6SmcDpLz
GYTn/ycJtPJ75t2fwQ6KQFqB0keZEBV8+a79N7oLR8DJMVuW69xopAX/pyFlbf0i
VDVk8nxZd6MiNArC+ejAz+Qxw41zOsOzTpA4TlxXZL5h5bxE90j25FyJud00Dlw8
bcDlLwuBe6GJMCY2d+Pbh19TCkHlQLzQ9zm25Ikd0aeLYBnb4B47UZOxwGvazHhT
dfjFEsQyLkHGP1Gx2pNl+boHpUa+Q8VKGDtE2iFhqRsoIRTY5BH+v2bL2lg8rmai
SS2fydttjkkkmH2NQZXA/jwtAYvZyHQVw1mxuZZjVorxTtsVe/dwj+e7DI35iXdD
YL7qZ9q9l5si1n6SNZvjtfqulbLSpViae1Xa+vhiTugcUNEJOdFdSQ2Qn2glb8io
aYQkaKDgZppp46/d67YLkyDj2QBgrq+6lZa6WjhU5pxtaOTXmFvtdprWT3DErvc2
wia8VebFd9zz95PcPTT7AGwRc9EJLD0ywu4SHwWN5auy3OreWJRsG43AHC7MLExA
dXS8zQ/M5rSwsanD+V93bjenH6CUobqQNs+TQlDc68FlSQ3bzaCcXvw8x1ggFcrX
dxImQZ1Mqbm4KMyeeC88XaH3P40q2wFA0yvhWbq1o5lhhRkEqx/WeRIIg6xjIqgz
pi2V9khIxcTlsCyM/f51+80Twrnl2BFm1q7UxXn65nxzXnuZKFo42HWWDKA1HQ41
r4Of6GM0Q75ln5lR2owuWrvljqAmQXvbOBLhBeCIPeIDPJ3MVfiC46WWO3Ztvtfh
7PHbeg0SiS3ZV415A/5yklVF5NyqskFhNxtdJF+/pn6cEp1wF4tAMncXWz8I7Y+E
MHhLXrW3XRbg6rzvrW2MnGJJWiKOp+f+6O+CLp8IoiO8XXApsvZLxKiOpgv2Hnbj
GdWIGFYhCwqJkmvsDnmrvgRbQ1rERdUxdNWPMklgauLpp2PhfWbHwXoVGzhAIWIF
utjXlbGTQHB4aNH7hmpU38OjsuW1Zh9o/48L5vM1ucIo9ozqy2d//wsf6HWxg5rw
wsbAFRQjCgoB7GnfyZ/8hbzhbqpKL/b+oYZr4p4WNKRdqs70OEPUn3aQVBRDs2Ah
cY27DwoqjTBqvI3SiuG2TOAG2mK0GUGjNKWVgf7Q7kqfHkWFPmOzp34J/qulTJ+x
6dqOnA+DH67S8BJFN9jXcwpkljvNh8erYBtGpjFFBISEt0xwaghV/neRbq1n5/dy
hcnXJpoUY+u9X8BO25wbvClVAITQ8Sag76+DUaSgKOCLgRiaer9YoVtbKTHg4XQI
BVUDb8Lt8DZQwFsaWoEzWJ68zMh88hdwiSK2SxlwkOuH8vnQcaFFPm7L9CaEHkhf
8MRle3HgWOzCu93JNKc9WvEM9rS2Vbzc3Zl5LmNPh609LJlS1cB7QNANiw11ZEEF
aCm1ptJ24YQFmHvreswpQ+Xa4kaZQShYlpmyqljsj7YinJtqhe7asj8zwP0EeRNx
mrhJKxmic0V3wt3absT+T6gPSNP2Eppqtv48udTnp9vXZaI1/YSbUW2rSd2i+62z
KG3Iu3w3np4DNG34ZMVpIchq34RZToeF0VdM865fmf+82ezTxtJcm4GLswJ46QPY
MH7Ccv6dDNzhQE0lDHWevfBCbqD6GdyrEhLn6lm+XG9BA45doIH4ZxOOUwNP3fAq
8U3DZrLgiRMwJ370COPfyQn2uvq0TyAtQTaMhSnzYnu2mjWKw4aMLfbvq7kNDGR0
Lcjt5OjwTQPkjGOriMsa9520qZ4cIW+NTIihyqqzTK2aN5vy5KKYN/NxcQVfNBui
/iLKbeU33oYs1V1ckfzSKONTHrrnEcOj2dWFktD5hN6nLwLJUXen+l7AgocEKtgW
bpJ9C0s9Fch5GC7C4p3CYc+uvHoSF61YzAzYNjmez744/58x+H/4nQKRvdt7FeqP
GdXZcFgtRynSWHN46BBaL4dEKC7IFMjgjnseoh6E+DKR48Fadat6FPb3envbG+h8
uE5a3/35TmL0fdlseaha7FQtfO0t82ldaDMlIC5X3RDIQLwAx1MHoS5Ytj7u5fnw
tcGtdeN4MK25IQ7EqqAQV4tXdpO1xfzJlMlx82510gQT33cxI/AUQajJMgd7CMjy
aDl3GT4tg+0VJhy0HpcT2mlX7twoTR+e9dzhGviPd5mRXB1/5NooKgFE14J5sZxf
klGRqWbxQdbhRzv4fedtZ7Imz/5+DbjlAJzHNV3Qhgzh2L+drXNOVI142ealKCZ8
A2RFz8oqgBXdeWI35mKZmkWElIVM0nTXaJTp7auzNsB4uxKcSMwDI1I/MAbu9FUd
3C/hFciDc8Jtf3RDyyxLnm7tbjyC2EKHbsdpUq3ygB3n1seD40ARgQcTICZ6J1Qr
n+iILM29clxluhVOHSatPcfJtRW1TB/497gBVs9aOQ0OuYg5sm5kpB1qcZQvdQpI
bDeQ2LSxszxF/+m+TvPO0+iM9Y2o8d31Yz8+uHiA1VwKMbjmcrdnXT39py5U0bL2
wjZaYtgsSJ/XSAZEl7dwE7NSU+R3cVbhtkXGcgX6o3/JE3RTlEDtkYSBm7lA5avw
cy4ENw0AodJMDnGqCR8GD3BBAcoPYRUey/fmamEluLAB1KUnX97aEnfXcB41QKA0
kKjKKK8iK0/MKtolzW7QEvLTN6kiJNLrbxMjHIMbwDupkrzScaPnANS+yH+jr5KQ
w0ln2v9RsBFkHu2K/mlHA/+QRUHskQU9D3m74y0R5Q2K2mG8Ix+8BvmAu2+Xzzh8
ElL3UTbXO9VU6goua6vGdgxte0lW+69Xcwrq0kX8orxb2TD6rz5qafGGw3p9MlJP
fu6zKuIU7YOUX9nFEm7VAE5a77XYqA0OZI4TzGoZ1DVUTDArzpCybEAcVVQIgaaI
rhvsiwuWFyp/ku+zWHHRQtdE8BIm0K4x0a01ITh5x1zVcEC0dlkq7srulGG1XD2/
GE1VdQMxk5JwMHel0cQTBuwHgbGqkiDN3jYYOWj4BClTIqYhpEHg2jn7DXOLw2/z
kL6jacoVmO7zwQXq+WMBYVQFocv1a5q2VJc/bbJBgQwpt+/mpg51VQ/95iYFLApY
36sbdlEWk5s3G4AR5eJLjL6WitAAwEi7oJ7M4ax2CTk85v7sviuPq5rGcoJIBusx
xadlUMNXRCGho6xkLXr/odYMidy112fJzTPHzNtHHhunO1rosmjw7tGRoufHklFr
3MY4n52XkIpq3UI7Mf2N1xreHmONK7LQ/OrC8yFj1jlUBtsEfmVUQEEAta6uc1UB
oRRH3tBtpAOnAunNFODVkCSPQFN08dYTuoFWeWmnpk784araaJXctrYdQO323g2W
8H+oDmd5b6v9PMoFi2LwrrHB3wbXmGV9ApvTMjG9sgxvB62j9Uoauh9JhqHg/JRQ
xpy0aj0XP+/W+BrljPeW62nCtcECeQfyKlVsL8XDipP7RvwFvy1Nn6bB8ez+SqrV
GVabg+G5Oqy/rUrGpRKVU3mloAnOAQU5DjYV6o5eVraYeSqJrEbPYf8iGDfXg4mh
erBJ+CNKRH0DLW+irC475hExQtflcTtLeq8LcBa3lsLcJRCbzfBuIG+y0o6kihaP
V3ZGoymyPrRDwl+zJedxv2zaiXsYREYZOl6cydddb6nEH9w+fAwQxNEEd+NK9xy1
zxiZwcgB+8BDij2dPUw2jUX7fVxHw73319fTB/NcjSdU+vNRK2t75gaclN76BI5w
0mQFIjNyQTeP8IWAPT0QgH+vhjDjdYtfZk1yuru/y+YZ+rd6LyMC/is7TQPjciul
Vw+IXcpQ30GX2kM/2GqXKfGz2tlJiPDqWQrIdkFjDwDwb6ZhSvT0n/b+irbXvpP+
orVbnaG27V4DVg/JraMhp4+Z6xXAQLX8r/oPq+k5Zu+gfB6Ecpo7rMROr4rUVyep
N0P7qBaPDTuOmskr06pwfOW+Eoc2sHM7Cl0PPd+FflyFbVa0+747gheBiu2/6pny
RJ4IzOt2UeNJZk3QWFNu9oivHeIHhyDKOA8fFQslJ7lgvW4hB6FBN6P2FX8y9icm
hlxOM0oAV0Bvi11XScTr+unWwyLxkzziDWxdVpG3C74iARhTiJqcgSpHEBDecXJ/
q/Nd66NgqBrG7Ng7JiLURvxYBOGtGsclUEgWyBs0Vv5TpxAFh/bl7m7s1GOuJs5K
GkcS+ro3drRSl0QihPHmKlodQ1azimtdQAmwrsYxpApXCM74uVnZ6Sbj8c0gWnxe
3017efl+kkLDA1fYaB+ZKtZok1l1p9sgUuCalbOMF9jRshVjf1R5UawRPszgsbcI
koHXTsVccaSrgJz9CVt0Y8yAScCh/ejqJvJqccJ6b4utu0eXyWY1xog71AwVA6XW
jAykzg28p0WkNZ/6aappjivVSQRlFQ1q1asJ/D6Yb++Bk5yJb1oUmdx63tl+PGwz
tLlDYEFYu2J5VIXjWg7C3f/J0i3YBvAITcFR+TsMMWOT1A+KpWwG0OBxSKwI/HYz
hTkyp3ehp8GKHOpuCGTGRKau3FpsqnFEwDY0ilMeTTMzrJHodRAVolxrfzn5bwTr
Txid8qrme1xD2zFWZ4mvSKFSh/dq8GD0woF7hX2jjEzlkP3/+HW2nZW+nKrg2spI
ib7t4F86uf9Gm4p3huVoRmMxGgUbmefV7a8yxKdfkDkDfNTEL+Y6o51sS29jRpw4
cugRTePBBrgRbuZH6mo6hMgxL+4JFrCIU5QH76yigtCbbbGLizcNd4uZPDD7HVD1
6XLC8sWc2Igab/JbIyJfl4OnBkP2sTGQ4laz0lul3/veojC6rb6uOn8RmOt9mMgP
UJDlr63xcgigH15T+exapdxS8kesZpo/Z73IVEAfcRCCobuHZlrN/8C09Lp0F8dt
mnV10sd+PW74NKuBAU7ko/f2DE0DNrlOOfkLBENVfTe/qwXaPAP7+qLm3py7Mmxc
olAGOS3DubnHzLjHQ1LJ+tkJiI23eurlf44DMjI/Qwwot7BlPXmtC4vsQ53RRwMh
GDMmy65QcTcuvKS30UzAttuD3fMnI68mmk1Ijigd+yj4IZ3qv3ZumyNbv9PNsG8Y
L5UT8bBzOSxJE75OUIVtHyM8jsr9EfeAEUQsuxDOjFITeYHL2JfjTrY10fqXj8JZ
33HWUWDov0DOI5fzhqOy4NxQI8A34An+5KmkLkmv6ejKnSCDQiOy85E8zWdRqpii
6OTz7rWR1AkGsgculkrMZ4TvfFWz0+MSqufbMsI90COL7qh1o4GTZ5WC6u2jnb7W
/dzJ1Y/8bYx3hKAodp617TCmZElPY2xJLk6hREYjcNgkLWy+L+mFCfW74I6PdeyU
QgUZ/xwKp9vtH4p7iOZqGztCAIw19mkAY995wBDrtbdlWur4qdKmGF1eYgBH7SOu
5GBF0LSPiI0q0S1dDYCiUk4o5LFgUcEArnm2sIQ5Rdj685NjIsneTnKu876ajEW5
FTZhPEWeK30E5ERP4S5SxH4qywffWv/Pm3rRrvh9u9LYAsXrSB73KDlIXhS7ZmIW
uwb754cPTL7Ikk/+TLMc0HQOdpAP/bc3AOGixvyd8nHyaLck1La3phIFhlzOcQSY
xtMtQXM/BFNoH/KkzZULwpaZ6nnViN2GVf90ZUrcnFekm+BP+5im9owGmHm0frrO
Ct85vqF0zGS3WUgX+suLkzYZxm5W/r89KpgX6NUq2SlT7wKtH7JDiUSg1YQehmbt
Z5prpoJ3HTYVy6ChyRB/Zf2cqRNnDkVng3LLuTf2YS2WgCwmrl/fysbbkeDIWKXt
5ZCBwuSkXvcP9aPPIiut4+Ko+pWBFtdYxRe9qvWJ3jR/ouzuACKxxJyUmRaIYMN4
AaP9gJMszWZ8jrGRWEQ8LoHR5Itx8b/e7jrjExPr56HxL3g9zjSKDcaLGLI4qFy3
sEo40MYtRTqZ4q1RmIQZwsnIJOWEx2Z4yaxoXf7ICseQCWVAs6Ig5g9weL0ZpUir
+zlTcPSQLqOhJEA7addPKICEKL1f9jUxzXBK+SmMqYtZgp+wD1UtL1/QJPGmjtfU
O6PaXVOzBDGeMJm3+WxScFlhAyv2+iMVavRRLyOOjjnfpiX5l/kwOSTmGPu4ZZB6
MVF51T9TMOVCGK7cPlDZmzwFooO/r3pGFSuM7WpYmRe4i0wIfNBDW0v8lNZZmsXB
CdO0r69WX+WENZXe6rlyx+VJj6iNGYvXI3wrqe6Ja7ZG3aOvB/rdcfO0R2SHNSq/
TP52CS571C/whjAtrd/JfkJttM/8PqJ4cdSfq/ZFhtRHzi6o09aPPDhZi0rDGau4
HkWfVhkn7pY9EdzIXb0EdBmK26vHAXYNMjAqglsQjryTFQyzr+gSoVe22KNsG/KD
CDYlflm+bF1TotLAKdtJd0c3/D7eHiTsBNl4/rLtEuethREqjlyI5JwFOn/5dSF2
uiBuUDdaKl0YmERgGr2sreMJQCIkYG9GX+CN/EsOyZqDgpvpBmdYIx5O/7HEeh6v
emM2NiiHicvoS5nE79VnnEbBBrpLrIwwaV9GODUfSa4Zg39/sl7rzcjrrGfBxmIn
cbr1OmgjlfEASI3Ki30HtNiqmga43L0IiBwqpKlje2URB8dv8TduTfWbeZskz7jB
qy/nAjZ5cEFJEvcgp7cOu/uVAWjphTpMNEpqV5MEBoLeh9ukm9BY9dyl+HoiZXWn
co4kgqpmcK3OsKrwQoxxbB5obhzWJN96c36n7UcLP+VBr0R2nB5Xtq8jL9CPmZ3N
zLwwPYQX3oD4Pj3YR2CvhMMm/X6XEYRLGvgg4NcsjYBNkgalb1UNbCsNk9shBjOW
1gjD6zfGXn3IodC1Gphdp11cpxJIxfPDr0uamVAdMUtaA2QoCYdOylKVcu8LHuNp
QblG53rUjnDi7tuhKvYUSphcA/O5B7MeXOy6d3ftcY0P8S4Mc8e2HY9LQic9M9ot
thvAVPSQoCHJlTxTmIePnrp0erbXtaa2gu323JGt3I4Iyamv4rGjxARSU/dpJ7TW
LwJKV9DaXNFCpaB0eRvYzZSswkmJCkGzzAT207D716OsmUW+2g0gytLLADBonKvj
RDnphNLbdyi4Z03iutmLkj8IG3UuWJgaiofWukFqiQztVdTRUywssnEE35yfCMWR
nKOLCbDWszD3ZWNg4862tyB0nrvOrLBCGVk3RSWt12xk6IQuqqgVby5PMlKyDOWG
H3zXu+Hkv7T2gg9vVmFEwAA3SHYJWpHhXNEl0Q0VfdO4klIBT9wh7oMnMwiVTw0u
4Eq+v3edXW97GkBTO00e79waYqAWXqee/15h2Fr7yFvX6z1NnUxtkxm+4WBlH7zm
0z728YUeZEm1A/Ogx6Hs8vmBS/ba67vNvmZFKj5WPzlplbM3kfaXnQGfDZghsivw
e09pK2rRTS8PzRJvsDMZWjTmsLWWSj7KmXVT00TdGYc1nN/OmDEt7jEIJmW0XReV
NuGDAkNEQOnqd4a+HPBa/YAud3R/3bhwqzFjpF5mDiYu4bSEss92d0paErUDdgw9
WylOG2o1umHOi4K3F+WYapXNo8EAum62YKcROfF2l80uhfntRllZsVqaJAZPK2Dd
8f/G1ZNZ/3XoCWSNjzhYpW+thE4abKvK1QnaZRj+HJ37UkDoZ2e692yfgNBmvMca
WGetiCUPqXFKxcysSRWLfnrTgRxWdOm+IE+W3AMszA1hR1LfshkyoFWCHBgsOdCI
Q+qcDdbjCm8sBsez01tE55PUsRUbf0y+FwbGfQxhhIZmilNRBF8GddwGmqLU/Deh
Q5aED7NEyIJml/GtINgh61sRSeMBCttlDY6LRmFNuA7mcwBnStUwgW1FoFUAl19Y
K2l61oS1RHC5jLLRWivRQ1TkwGpLdDX3INUMSoy8ghMiKURBJgG5bsSqu1XSGYb6
+EfAFQyi9oJ8hVCuH/wbGHhwTVRNPHH3uNGdw6YnrUACt5gg4ZXXx4tEeXgDR9Fy
0aXqe1Z5yO25yWC7SmvKkqLAYCDsrf9rOnMdDZ7mz7VCH/ObZfZLedvV1U7b+VWo
UnZZS2Q2UFzn9zWqbm33IfIrljjR9Yt2o/n2++7lRar/zpTI3AaBogYOfIvI4LPk
6TnlSRQas9x3kVpCF7OWL5SwIzolwu0SSdEkteRym+AzV6VKsMHakIZKC6Kkj9m8
xdNe6X+0M95ysX9wX7YHBItNvL2IEmiJs1IB9eeKQ1noUcoZKW1ohvtDMIQ+gvaP
3Gwf9AAMVj04Oekshlv5M2d5hckh8efInqEkNpFvQCkHTEqrt71t37elEzP9Gd/V
NTvuF0iQUkxXA7eEZRK+8fS8bVRs5GRI3qVGZ9JI2NoOYiW4GQ26IwlIYt/fhZGG
zgK+z844wYfqZOY2WaRBBkd7+OHJl6W9K60klPLROPEJCtvh7BqRKAAp336cb3PP
+P7TelnoaSLEFGm7Yxzq7iOEbgtLy7dOHAAeYkU4o5F7SgRlWGUORt4uv9ainnas
gqkt108LJTU7hroM16kIjqyMeSR9cf2RSrh7DeI4ufX5wbgvYIKQWfHL8ufTsWog
zxfX47cD9g96Ho0s+P71qCokqGd+mwRzuAflYHvGwqoUAtQh5w1z5HyZLr6kDrqg
78HFun4g38BMoAG9n79l1y3yaGktvKP9sucKMXSU6xSwNNVm6JYLQFXWrVWBihc6
5EIXI6vrQjCqtO8vlAhWIsMICywpO917IX+IhOGOwflJVxPca147C7rtyTFXVJkx
dor4KDszomchEbniCyfqpOIz8u00cSZrQjowOAE6Ver9B4fXBRBI9zjJTeX7YEQU
Vz5X3/dRzO8CoPQnaNjUAEd/lQDy3g5rF9NGqpD5oWMTb8SMRRig7fpfXIcV0n6T
l/vGPZ8ioZM3LmLkWgEJlYVgaY9xpCpW6XggoEQ2iMTPgTPhjrlKw1qwldRdgRi9
Rwd2FAzVlEGa/jt7TL8IMoBjquZb3wICpXECvMFFgw9ibdGmm4oIgoNgh2Htppky
w28x6ImnA/9SRjWdpkCI4xiEdOGrUPp75gJkAtnZ8VaD21Tpl53y3+IJCK0ons+W
16kSAZVrHmUfG+b4hjjz73+NGvrmd/hMiE2uO2zxfLHdEZGWpwnjuRR8vodNRUDb
bgAx3UbaZHmAaKIZpV4SHLg68N/A1ra1ex+sC2cqqQ8NxZ9JP0K3Qpx73xu64KDA
7Zs54hpdQveEnvbiAJsSGnVipVxcOmcuaY7MnMT166l6yZur64ER293ITFFMJlX5
J8JG8JCvWN18oQIMmOB4CoF5fZ9uIxOqnAngKaFEHNw1yQJ+1rpR+0KrTs0DRMIK
5HRUGVaWkAb2rfBqcy2zCsfbaKEtxvL6ODnJUKXQhLkcxAWJZHx/MqSEGXNap5jL
7MbinSu0+WF9IWKXxEqDKzFDNFp+dvX4ddU6vecZuAEXQAxa/3435Ff3jb9D54jb
ErfegsKSYDxy+eXGfnSC8SihC+g2qk5j0ZCfJW6uzXeYcGBBAefXfCh2/s0ZjtcC
m3kff0fZDhSWrQQc/vQv+FzQkM89JXmaPBzpU0n5W4x8E8Kpv+0xBa1Q6iMlY4WB
+w584RyIklGGlmSaGdpNAod60dKW4mUuaGgvNURq/MTKdt3cnQvzAAgFfVY+RgxI
k/Ych95P9WNP2GKVwUfMk0WWcsW4kh6ptwU7F4AdzZSOgWHB9M8aryybEb0Oz0Bp
hm1IclpbezlmRkc7h8nGDzg/Tew7zyJQHarv+Mkaq/Q1hyzpw7fIoVWn2kKxSBpy
VSXhF9yiPjwUETEXHp6CYz0F/+jVFJAF08esSmT2RyCa5afBdnCnHF6NiZPRrf1p
drCnEiKW3lw2cq68D1jX+IUHlH+VJru7fWEIIFkqbpLdKtJDhKGcebUW5GeybXqo
in34HI4gSUO5ZztDhPDieuzBDxrbQmgqnkSAoAYN/E4fK+OFVueYqrol6W0bZjR7
BPqcCSRFj+5+jl9nxX3p56ed1MKCk4qO9MpB4NRpzrR8y92xEZwfWD1tF0Ba7j83
7f8s0r43bccIutQnuAaJiIXB8mCqaHOZ8FT2fHAz2s85VFmDGBRg8cgOtrK9762/
zJvqtCd3+Cy+SwQ+ZSPbmzHeSLPjUani9HJ5MiZYdJYF62SsvrAq+QlsnxzirCuJ
upnWUhdJZ2BqAEqxtchRqKxY1u7pjADaI3hBpu8RKZZYw26Ak1VU40T5e1akBito
mtFK+zDrqWnpfcs1iZahJ3nPy92G5E211990QKPnvwRw47Bse/bnTwIbFAAQnmVV
yzwisUK2925VY4eF1M1VedD9airI4mciuLR7ihgeybl/GMlRqTOtK0RhK8FdNxaF
f5j4DHvuy5ZrMVCd3oQWEM0d1+AGNd5XBf2Kw1ba20Ip3qZs8L2zI8YiMqLflJv6
3CNcrc2gIvB5TOYWs+f7KCQR2qmbmICkTR3s4RSI8z6gWjBMXUOKDhmdoBv1qFJ4
sEZoGjgZU6IUxmpLquVCCoKOBYqwUzGKBku/y8wmK2xHEH/xLj9Qp/jDBTMdcAFu
3uzuF4rppKxuUFU+zIJlWmIohK8Arf5PSCeacEeIRHubVFsIWVATnWj16kjGZqDF
KPPLJVeBDLC8eS1Kro1MA+Me3NF4TyOmXYzG/jUpTgFOMu6M9kIuOMR6HKPhDaBI
yPDlpP49hR7QRH00Uygdu4md9icLz9suDA+KcVa+zDrVoCduEm5bb/ZnAsxPOogg
NSj8UzHhpRyAKm+PxD6M4LIaSYRXGcSaZXFj/i+mK8il/PuTkapjEkof4T0qspxr
z8FoQvKus7V8puzXzMrkac1zfTlTX90FWWJUgN196Sdpb8z7kvyNOt2sDOEEybyz
6+JO5BAo8pHN+xHJjYTS6as1OXGQt4cpsVab85M79IpcWPLDcggz1jXj2VUJL8Oa
w3cUbqD2Tef7msXLsHDRrkJgwh/Jxm3dXg0rr87qQOl2u+DKO+DiT1PG/be02i77
/kbDjM3J670TOC3V4WlYUGmM7LLJn2gp2dE0DIgrB6E3XTIPJR0OKTbs0L/DYjzB
4ZePKLMXL+Cz2rkpUO4BpoFpJ4iupX0hoTjEoEtNVJ23hJerogawzmKlRGFp3bVM
wXfxi6hdqoFzlTL/HmVTuJZLre2OBMce6CHu5EB7fUBsEfpSo20BDpHNJKssr1zP
3h+p9ZEIbUmCf4ZVH9sRlwGRLiFREnShjKZeuMsB/Y/E2a0ry+/a0VcpKtDuEHEm
ou6tiCX6LFK6oa5NkwOxTemJELJPXGwYk3RpNiQ7VA+Vr0fI0o34P0OZBBOTIhc8
EFtottwcLsat+IHwIpX+qi3ENCn15ehs3cPwNt+sbPU9qaEKN93D1kAbWG/VLa5T
qPZJHcVWuI4IVlwTPk3juZ4RqtIaAIJDGOULCN3wwdfZZf4WH5GVq4Mb+/+ZzWuq
cvJhXY406uWCK0wyROJswII0wKinm7IwwvjrFcd0TDpZ7Nse6xUpbA1wqAS45QPo
E55wRC7boGaLUWvbs3GgBYHDf2MGs8WSdQBAx4PquKYOPErEjcMaX7cvGZPCjk6V
yVHW57XijNLXCEjgdVORSuGpI5fiT3UUY8Ff3xsDZCPleNTnpnE8JKfU7pxyAnh5
goXV7x91IC4RH4RtBHE7o+IdxQ+RUbzAMT/JCnGVMA997zoCvZPXwMNoLzfy0VnS
tS3DkxYG1IUA41cmADKxjqDtIqktXUnbf5AoUwB6HSyaI/5DBITLJ+nGM26gbaQG
+X5DBofRb3r6x2I5prHG0t5nBYI4VrSPHYI6D0OOPzL5bcy5+11IwuTz+XhIxdf5
f8dOA3FqeUOXHYRgHiv/9lwFzhsQyAD4SPThfRnb0R7JNNPHa5sFgbMWpSodMJ0g
iDf7tKX2WxVxz5ktUvRHIrtnbF4rBOibPp9Fucu+yq0vPU667+MX6Si2XDIKpRHg
R2+hko1xHxDTT+hRPqLf1OOd0Xd3HVOfL2TDSS2WnD6NWsUHIQcFODx5bD2ODpJT
d+g8VOjRyYxFaW5S1IcV+SsStvX+ngC90Bo3DIR96qk7bEmKazd2sgEPsh5NqtBj
Kqf4Vp2pIUj/hASCd+EyCbybjc42EAxxHGjbinfDOIv7WwpQ66wdU2Xbp/eJ7XMp
a4CBI5trPrfXZ/sW+enkO15Rg+4QXbjXdAI1GI695FBO3CmkZ3KgGDowzbM9dxJ1
ukIc7fgR5kMQk0zlcQujg83+UGlY5qloJ1KvyLaPhvSGRvTP5tZ9vhqEEoPzbD5i
vy6UnulcWGt4tSRCYbqo6JZbtmO/JBNT4ZjSij4v/EdOizn8HIRKyWpwgrDXtEkD
AMgO9l3JF/igeoPrCqbyVBBhFU9xVNLBXwHRqcVdvH7NfUAO+hN3VCuoeD3Fj/5I
KdgG8ZdTdNMFnztVkPAQArpXmwf1JV/egSYk2AEemDU9MQ9piRlDvp659aEjZCrU
MZjd+xitnkPbfQ4Ic5IgK9KUS9/76XbEhD4SWnjXqmg5QNro9ZkTRIHGhXJHxAed
DcfYuX1jdlF7KyE/e2YzOFwC0yckdTV7D1v/7VWcFtPvB/DEkOelIA+94rqiudys
fezAFpRhjodjVb9yWAOqyYVhdELKuxNSk1KDQDv4/0qK6C6gHS/GqCceo6GpNNDc
BhOFcDlCNTpsGC1xvF1OFBbrpcup5HQV8ok/sjOXuI4sjPKkycCGRyRkH7sHpxwS
n7Smw9uivGkoBS2Gju6BWBYrXe7nwsswKnruJ+zcZ905zj1zOsthCfBvintDq8JP
LEAXUFCWGicp3maIfSi9+6sNUFXMInFyt6ekNNM8Ox+tKXJeBI9qa4hB2+raSyIr
I3M14SdZwK1SL9Uwi9HN8yLen8V1SKKCb1wPl1w4noXQyjnVBsuSAaRzFIbdmsLB
MtBOfYBHOtNY9cfuYRoxj/k0fX52cQr3xBG0mIFnrRU1Y7CFBdJOQ+n3XcbE5IkX
bf56Hdh0EpFKCqhuUwJ627jqEjbtwH6mEnmzOxuO7QtxuDGevKGjo5IgeoQm9pC9
Z3d41IQTmKDNkP3b7sV/ttpyOSI3GBGSdvwz2nnn2KZM+MkJ6VEYg7x27GwzyMSt
5QyBvnE3IcR2tcnfZ0CvAh/MO9dWwaLdguwxPCJI5xbfVs3JsiCoFGdT1m+pwL+l
jF/Z/j97v+EM3VHA8qcxaW8VIJZF/iZ/i2o+jAret3NAlbAqG0cWPYvb/EIcbsCz
AIjVX++9GBwaVfB4yCSjuA+LMBlr3bscY9zdbfXlkNbaKQGv4Wm5ahfWnsMe2FAs
gFeK8WFc8aab7UM2x40Z6eftEhVoj8Vn4ia6aOZwo5d+peixuzqiIM7iOJxdKPt0
XDhGn2GNAFvInyal1tDaf2z4GX2mb5+5gcfuweCoFHmE35m3WgxSCQbjEl4+N3jP
cfNy5PiW3sqSJ+luzVgLDl2Q02d6PIUpeNNlJRA1FWbSInP1uyeRLJK2zpnkHH0T
/ca41gjpY3oeDNPGY8aC6axotS5iqhDdk41i6HnWSmxV7sxs6cUabZo/COQ1gIDF
8WZzpS0qo44nw4kKq4rToq6sKRR2xdyeP0lGf9DjXcL9ekwDG1jR44M2mSwtVvhH
P6uaPa1xr8hqMvWH8OCpfmePdVExLu1L5LWmmwRsyCItj/8wuNiTrhoXKCD8Sxq4
KxqU7IH6gwmH3PzwGG7dVrkGWWlfmzweW42bslFPuRxDNi/wGlNeRkLOFnboeWFh
f9I9LNzRrKlFs5S/dSxYnNhKr7pnPgTzyqkXKL1x9QY0+APAdRLQQJyQfgxJXttW
+NXqnq51WJPMi9VPSTv037DolM8p7tL0Pw4UrV5vW5i2xjSBArRvjrbwaWJNYgFV
Szn9OAYQkuzJSf1iNcdECSqNZVpC3LgItxzIbPI9XgX4x4HTxd044dEodek+ow2t
17zWWUzJlIlEyOC3bVVAdwLYG9Y4OtH0LEQerE/rPIO4yZaiEgFYxWHyOCNaO8jm
/pELPA/+rYJfxywrH5s8MNL4ofBmruQt2NQntahD8rDBrIV4nDOTcYckv/3TdIV/
/9p1SnS67C0zoC1WQybo25i4x25+18vrl9VlwyYgUW1DTO2Bc34cs+l0f6L1nBSo
aTaOkXeak4DesP8p9uGRx9hwfe/mH5WD0yVQNQxvqjXIaX51vEqttUMUJZsiAgjj
HUpZN1jxUbutvSeFvA51xkb3J6iqzE4CKlN1Hxlce/AJho/V6o4XbyE+DTGzgXx3
VuArTRpowNX8dh48rpsePA==
`pragma protect end_protected
