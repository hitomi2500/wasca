// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Aalgc6dNDhbbA+5Qo5IS9UoQtXFrhh9Zh2m8YdcLunMa44nyji5/Mr7PwyGbis12OtQw0t+maiiV
pdHf4u4hBuonAdKPhlk7mPaKz+VD3eVUI9S7JG6gnyOIRy5zmjgiOjU7/x9A9ZmbognhySNmwkHS
k7/8dibO60+5k/LX6fH3tdKxT6XfnXxUIe16JPmJ0BYazTLT/GPod1SDNXFTPW8yXlVsloEmkT/D
X4A3LN9EntE5S5jpC+asSS79Tb+JK2BndAZodEHUVB5wW1089/21v/JlUwMZLxsR1oKWfcI9b3nz
8KRRyRZcJfr1EWkAKXxHjfdtqRokXSGsen6m0Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YhWpJwpQM5sNfOJfEtAU0j0Ne3z7pSyKvRcoOeTNbNT0dioLZGKpFr5/sPA7xMA5jZwa74DLjO1E
2URWcCnt2a4F8C7uEaDRUxCvRF56isZ/ySD5fjWjGL0JB4EXqwDypVC8grKZtcjidZizT0hbqnvH
IIMGsrUzmzM3ta9WOjHEKXvSdeulkVBs7+NSp8qdKdaa1QiA2T+2IGd9wVMoJoDGv2Fq4XsnjWeB
VaPIzXX9/lXwVAAir4rNS81ZOR6GjZgOhsS+IKAcgj+zjMuAgS4gfbjWTDp018Wa6wrx+xsDpd5X
wM90vcCioNd1Tg/fJxSCMGAHnL6K8PjNME/gT7ZjPqf1BalmtLswfoN/fj19GWtqspx7nBnBecMU
jGaHH9mqIKkZ7LNE+CXzIUIryJxVkRXY3Smygs7kNlvinJtuYEpzrDnKCH0s/5wjaA5vT6PJJUyS
N11bsj9pDF4NHOQkJ1BU9QSoMKZMcCytuOuBpFbxuj405bTVFMW3hytRNOzUE/GimOTQ6TjIkda6
c3jS0+lWOq4Qs+FWUwiFWNRRfGJLewbiClftgAPx2PBm2Ze2MP7d6QNUkbpB0XZdnQo46olTbZnO
eH5QPwuNU0r3DgJd9CDfEfmgNuh8eLUxQkVvzLH57YvodetkfT+qCw28cwwMtfQhNVSrWPlo6qTl
MYFHQBL/WONaFs/FopkBeS0aPp+M24wRhZH6VJWp+8HVp+5GmXi2Q8Krg56xWTJdpeOX4lgfTVjI
6/IXgeZ4pyiAGty3XcFeWjSfr0Vt2MIC7qWGTODsQ4rhVZ80TXKmWM6xAK4b3oNCEeU29UxwB9sq
4H9cPUZSWjHgq2N/KpyI5w5gXFNuTEwDxv0F6BUSqkTlnltfAlpH0c2wICklPM+8N7Zmfd2F/djV
EFWAyWnXsgejljIKkxRpOW5F2/nfk6Q6B8K5JDnjTZjwixnkl5SlD5RXE7GhtmfofOfsQKDmqPXd
Gq6AP987sEPEkE496EBNXiSUaer3qGRLwrnYTY7u04S/8Fn+D1GjfqQQT69Q0rtzh8al/C1/Bxkm
+WofBYzn6M0/JqQl/avJTSws8j4cPH+HiFAFnhOVQa4PtnpfaT08H7UEXws3uXqZlBOwOmo6ofVK
zUU30gQhxspX7EC8tuo9i6TftKWekkctPKNZT/hZ2IKbdK8lOcmvF+QtX2csHdCJ7++s9UiJg+Fu
IKTKQVDdjdH/8+UkEYnNCukbIrKYJmZ4YVQLjbKRb09AQtq/hXyL4g4NiH9wwEJcFLVm+WWvFLZ7
NXxWjM1jkJU3FTd1UXSbuzyABju17fn6eS+rAfM7Tn5/BMraObO07PAOQg+VBnel6LIkCVn17GZe
VOEuuVB2UgNa9JpCaRUCq5p7oTtBzQnSn5ch7B+N3uP+0tf2GgnFfXr+8vsq2jdiYZjR2kKh5qO/
wKNADXvjIGDgt4UCHCXchd8to9rBAgH6NJH4X9m6UYUC94b+DgH54HNeG3uJFTtqyWXgGTdvC2Ve
U+Qii1dH3CKrOWb/r4q1OwlyvG776BeGZepLqPQI0aMMdlFXZfGMk20r+LsfcdffkRyo/mfAjmlB
FWWl0yMEZH83EbgM3S7kThono0C+sbS/RN0Kf1HWz3x++XJpaGT/AOhDy0lRL4eoU+AO8FG4Aq14
yYmVDRvSsrkK2QBCOcDTKDVSUKK0PFLiqAXZLBR1ewaMc5Ulg0ZVSzkDtSOxVP5H+Xy6MMJHM4bz
NBTa+Pu3Nmb7r5eNPhHCAMriUJQqTJTyi4iGwHjMO3tRrLmJ4dWcYek1NDchj/jcy48+CnUhz4dX
tdxf4TRORWCctUKNM1NzyQrKhCi6X2zucRcX3xrCn07V5YUwE40AAA4P3TRzWu/p5na5zpQ8naRj
g1Kldw74mnLAOhPAO4GaJFBSaPN3RCoNDWY1xqHewEW8aVHxnr9APM/BlpvnYo25zir+ObCxle0w
dLlCqrizhQPoi+zaPHFGt9rTUH9TQYjE4JEX40xzxdDri5O9mNvSfBWUyk/YO58HamOzmtDl5Qz+
DKae8+Q28zWIHG0UgQt2CNbsYRojpxPOErS4NUsmPionK2J+7vEYD/suc1hGxbIUxzizvmM0lOKx
Fa/nrNCiTw7Cy596LjbUAr/58TA5DsCPa9bNAcKu2w2R5WHPuQIuMJst18zayfuPdI8m+z/6Eqlg
p17mHMX+NXNip1ubS/Tr+3aRSRQo2JWUrhHMz3JsK1GGZh65KLnkbwUQPe6yHuHhyDeOVBoIgUF9
5IxVmiCRQkMZ3+iWoRv7URL1ng6VmbFw+cnrELLZT2PChz59GpIn39sB53OAkTmcY8de5JwVdowR
o4mQeCtI7Q9MqKb8Eu52LJq67ZE+hNycSm+nUczXgzlHlPhcnaAFYXO8Vw2/ZGnyIiRWBBhJ4gPo
9QXMA32DqhGfcGFpNE0+uh6H1Vxf5+7Pc9t6OcuIE08xzkWLn6828z7YKtMEtUlmzcwsjywXUsCh
kesJiCVDfSRNT8Oh62sNNT2zQf2XI5Z3ZOemHbQne5ms9JnOqiwWysoYfHPCbwcscwZK9mquMkOi
LHadOUInOuyz18HgL7mIoiZMDkQjO7Z/i7cltyKXXi9p2rQNnd8Hb99gNp1bf7Dc/g38k4epxaA2
txTrDwCwu12H6iSCrN48nUhYsMYrH1XKtNHBf+6XNkgaGz9dvKobpa3pVfS0wFsPHRL8E0uzcqNN
ETeXTKwnQXrFXKh3WbGyOXONwruLcTJ9ysxgG6cijeDuHRMOPtxnzsm0twTtd6ylYUDn6fZdv7po
lOLHEOkmjcyQ3c9kNP3RzwqlwTihxdOVnNrfNaudt1P+US34MmSco++rxdljHmHJ/8+T+dYiV1UN
fw6W+3LxXma0gLQvoNaBqvrqPpe3qVtpyh8yKRjEc4yi8aZJXSeuIQQJyrSLT2eUQZQu/SoG0tn5
AH4hT39cmwRw76jjhQ5UNcps3tEqoLqWs01Bl3BuBg6RoHENPojJlFE8MD79QOc3deqep0t1kgOb
Gmw6Q0hR4H5H98wGWKp3veqkq/nuaUEE9cylwiJ762krIRJZPfoB3w7Mwhn0PAssmT1t2a5ORjLW
3dXZZcJtinH2ZhLYwELM8NXnoHAzxZ2AjZ5pEHV0trKCVBHnBy6yBKAO7DcosFr2U54rZcqs95YY
rWleTdRqrmpJ5UQvxGDyar7SR3SKlv5X/L2UVakjaV7XkAzX3i0Q+s7znW99p0pLnxAtpUQcMqR9
nqBIBWYYBJYerZk21U17xDaTZ3Oxh0RLH0nWQJmHXRbpCD6y+Fv6/SvkrbK4XzuLk7AVGY9OHhPe
Kt34H9aalPNJGfg0BfZj0VrySWfDdIXQmCoJZusgkJQoutfJzSVnb28OR81bqU9hlGZHPAvkefXN
4zUrn/whYuYAV6dCRwyOf2n25ukAMQ2ngUz2HcKTSekNQtQnEYgJvrQjGaXfw5RyJqYwktqbnIWO
mFREbjy8/3cu4njiB/YSb6Zq7V5coGdTxaGvgbLqOQcclHxDpOQFDRLmouW+0qdYDwo4MsyQr82T
CSrWooomcOVVHbC9eD4DpL7SJc+ONGFyefb/jzi7tmNY2XE3v7nZ6UEsL7e2CYKKI9Rh7qe6v8h3
oBCq53WJuACEe96tBM3Ig4MD8w6Cx9SB16H+rWgHd2bZ1Vps6hL+IRtIVt0fkBkFVCkLAcpArM9r
3cxwpbS8mnJfKQz2X7drb8EiCzCt341oufxzxTeJiyiu59ZSktkm4pKWDMUcx6viCAshfMYD6qe2
X1s92CyAE8solH1Qz9Baht9GeLBsYxJe85FXfYt/THa9cpG4wGXLTYZ6jz+3cynG9BKxezDwYHVi
xR82BC7YdI4HA7kC5xacs0hZhlPEDhv/YB/+LveGaidCs7lHBc/IscZJGh9IWXnfh18rA5nZL+uO
LNpUu33ioSg4nYCxGP301VaQE/VFGW4WKhfxw6NlUxybV0q7Mt1pRL/FlrZViNvD1cwuI1CZy5ap
fVoeYa08QO3dAlANRLLrEtpYvWjvPLIDbRgpbZiIT8ExOsqq9t5ucV++HQGF84/jyAalJDoWcH9S
/e421jaCMOdiwpFg+5LRLFq/3i1q78U/WmNXIHMfrjrXBI18ApgDlf0/cfYbgDlETIgH7ANxn8gI
8Jsg4/vLcV6mGyVA+2AlBjzHlCWYPn0w3VUVhnlz2U4Q1HD5bzMN25zfNyAbKBJzfxonPspXMD+z
+nDldiOMQni7blBHKNy9GdyHzKHtg7ZDy0EFB3D5ygBtz3SA5XbOhXib3gZY/Z2UH5R/frLwf510
95WynYD9bxOfBJ+hElkk0yZ9Fn1PW9Q2gETX4ON3Dw1/7l6YeRBKs1+pCNg+3veHf6UBlLSxpzGS
foLc2ePnMolriEHkKS9PAk6GbQFNhW7ajXMdxL29N11k8gHrZlQg6AO6OWY6IKLFm+Dh/e/IMe4S
O9OOZOVlyT08YCTC3BQcCkhzc1a3EMXlyN0E32+usTE+QN61ahOM5yqoHmOjMz0fV/HruVGPL0Fv
qOwq40a2YfrHAAfmdT3AaPBzbb1cA7a/uiTwq24IpIHad6YU4w/2Gj6WQYu1lb57JXbF7BHSefjz
8MXNO6bXRXjA0+O5K4g31S1acSXvScpChxtxmlyV2fbpu/ButFjyLPKPj6Di5gjGMhhGADdV3DBh
DMhekW1wahl+Bwv92MPRD+rFOLaSA5XaIkoTXW9YikcMpTpYVzJSKVix3o2yCOB47N6V05zKRqGm
L6vOzKQEXb47oyAKsm+bbGuKKxNu5ZrBnvHb24nzmP48c4F9mG2brlJNLJaMI65IKwiL5SwbPf6r
GMvA6m2weqCI9pasv5q+jLQ1vug2sQmJWSfL2ytoqZ3gxJHCO/uw7aW6FNNBxbIGDQz6z5KkgImU
3JajrCirrYB30VrQN3SDHLkAnhqT5ysnRuHpDMKCLHzR4gr/KqhOE4DiLAMXgv7DNiq8YSgJxVaz
iF+z5T1GQmRkiJyhF68S5LqR8Zv+w7eC/vJqtGq58sZ4qXVE6oGGRMHuNYl3FpN5QFFvywKeTe/3
c1cGnmoFn972XVTm/N5ESUXCqKXZDReiotP74URy/GmcIeMBPCUle3zQwPUl6Di5UMLgZ/jVV1MR
rx5Sqsxhx3rLKnBzBn+KCS9bXCVGrZjNyLlQ9mLbxHezHpY5crbl+XaoV7OnNrS+pGZkjOK++Bmv
QZdJOgj7bZeyRu4f/Dmh+jTELna4XinYVm6D0JNwz8hamlk3E6Okuy+lMkdps7lmgXWy7T1/DSJd
mfnITggyj4DitaTxqfnnGM/1MFOhlj25T3evLG9R1c4tuCJA3fNxpMA2uwwMSrdBp3uDKQ1NjjnR
DQveCQo2E12OjmerjTZX/kjvxqugp4k96SDyeY3ek4oq2/mdxx8PP1pIBHFq9wstf28jN6SEgaDM
H9F0mJRQ8YX7zyxSTin6NayxUzbHY89Oh8NFAcg2G3CoYlgw/El/ybn1mn/Dze263Th5gsIjNhXj
ZUjO5bC2DZ47E0H1FX5RxswGbacfXFEiY20FC7zgDlsJaw4HaqY7L4Bm+swcyqKqVRVJsg9YmYQo
z37SOsRNV+Txr+4pi0mnw9n5UncfGrOnrh9r02+TostiCGSqVw9EMqveWX2kJ8s+26jf2E2Pckv2
a5UlmiS/G/2oaxf7oVvsYZtVmTsokz90bbmmOWns/zlQSoSL4frB9Tvu37joM3wHuqMSrCRKrF++
V1tlHwFsV7P58hwZ0XxoExlYEHoNYnVE1QDhc+KcEHvsc5KpMkFJ1Lc/n6c1EeLft7M4a3nifuIy
fUaRgcFQunVEzL43dH4qeFs9eZrGFoxKzBO2ft/8CayoeQuILvQrB2IlLo3q2P9IkJK6L3AQXBis
JieDUSoL3sWl3jNkroJj5J6asjN1J9BxJjGOa2CFZnc9v3u3GQLTFS6zFkD9ihdAzWnPl7xzojit
48mqoKsCkrPs3EQ/xhM6qFH0P0tHGZZXK1sAWYWt0E+FlRDUWMAlrZCcq+G+stex9gijim9ez7WW
Nqgcscr6myOhC1n+7NjcM0ZssgqejrDn7omTtvK9JwpQv98No8b40uObp+FsYs0OVKMw4yDlkPM2
IS99ZjCIcbPi7N3drfWMs1eCt+j53/JVEUePkpMyZL0/MFTXfLrCjiq7dlCxFFvYnn0cwJIbszqJ
UDZwmSqG902jdovG63xAoVaz1zdWJbAUKjhwhJxwW7WVLtB7SkwvSMpYIluRXqDov2QIBrdpx2Az
wztspVcz37iS4GjXW4MMD4ZCMhzJlOH/H8ZZx0oxkNZKuNtNjqfiqZmrIpPi3W6nvq+3g2+HPJ5A
yPsYHPrN5GVPRppdYCLvB+7nc1omWy3zjSBv0nGy2PyQcsfymvAI74FWWd5XUnwJYbxN4LMNr2tT
wtpvHLslzcqlMBIa/FuG5Ce+k7LLaFCE08Lkcmv9Jv9lTdptC5qD6eYOARiJE4by1PokQx6ZQfM1
au5TZ2/9l8dnMcj6b2qDwalBzkU/B1Ce9UAeFBVaueeyfFTLikQUzPXHlXnqMKXEyt+TgVIrKhrd
wYdgPUxI1CsYsOwqoiJneEuzSrni89/upqV8VPPT7JfVx3qI1zP00d6jK2rud7jPm9KK7de66YIq
6jfyjfaVJn50yjyCPUcvkv4/uSyuWWMXXkBF/BI6+75Iuw+wGJLsaMH2Q2Zr1nO2Ly0MBe4n+xMr
H4wazoZX+cptO+VeZrx37Fd/jmURr6IFtQpV7PAZfBlJ1/aV8x2yyGh3NxnXaxBXmeA/QyFYoG0t
5CvLfsOZAgLw/8pEr1N+o7D3E5KiAXJbJkkiY4iiVa/oCkeR9Tazb/PyBK0Bi5Gk+WPnnohX32C2
CstKIAWAefAR4P7I6we2vr4S3Eq3K26CRj2VioNrhJEAiYhfW0qHjB7PrdTdS+R/HEjYFzh4xlFJ
Tv+wMZ8SGV8pgQwQIGQ8l5f1HhhyaD2gidIExygsLnEzivTy0PeBxqRAYiJ2As0NeR0VMm1DbVpI
Qe25oOql3fukx/agEXyLBg8GaSpWALRWMrPgN+IMoMd77p64s4s+mS522ySDv/gFAoG6jst/WjGT
QDua/OPg0MBKCrunjZSLy7EbUeiHm1JxXoj3sCHKac7mFHhR7NiKqXqhbWOTRmra/ppJj827VBRW
QGE2Eh2KkRCFyalNAPqQ86ym53i1lOFB5ymIaYXnypBNjMNI1fBS+Juq/wWtVWOXxEjpS//wkSqU
YVi9yVJQuS5S8AuPZQdtdCXYlVsVwMYXulnqa4h3gpiTgRI+ySXDqV7LLG83mfA4aGJFlJja2jAn
mnlFPqxMta94FqCNW3kTEbkCCKEGp8FqxaU8oaLAwHRfzowGTdezBIhLPxPEc3ZN9wQQWHjgqDmt
LvbuLYyPPSDwcWPpgb+4kWyF2MRgefDnMNmj14h9WE4lFwNzuuWJVwFFKX5fV4PxLYiuTU2udp5j
Z14XuNLyIS7HdC1NKsTqzAuHtD5nqB4noGVvfopjhKXbqfvAr/T4wNKZuPdm9gVIrjS8fx8m+e3l
o0kX3oQ5+XAfFnaGGnvwDFxtA1C2VmiSIH8vxHr4xT50AZnpvVba2xrymjXoo+Gv2UVxxizXk11d
ZvbCF1C8MUaLK0RmCjsxqlXfWGmFkDT7rRMv/60s9SUqfh0Y2I3WaNYRbqGIaKlFpCGawRVyAzFg
PEb3NfzdraKYhnQ52lXfpPqtvxI6NjciasfnB9IHJ+bVxVU2YtoPVofP/rRFdokohQQP3gzJCfpA
CO7WNRjynzCiZJHLz0+GcGiR++ViV01oeyuznvOwLaf07Sb7OCVWRNBAzjb2xvbbtS/1iMzzUwuh
/nhBlhq5kv8v1feJp9i/T7sIDO2UC0K866xaLahU6BPCfdUgt5a7MnshVTwIyEUt906Q8JPmkMY/
NIv0+CkSrz0DStYgH6uPgKrQ9UOgDrT7Uws9N3NLwsdyOJ4VgBCVE2V7h9HYUJUfupBtFgtSry7S
q/B5l77ELmQ3zwuKxs709xVp65qcVDC8L9VwhEKrjzzYPZHD9v8so52QeZ59WUcsxIV+B4F1ahd/
xJ028sEJR7EvNyF+YFrlcMVJsTYFnSZjUfqf2g949sZe4kmcEbF0j3GsuGuiu4G+BTOhACOSohRu
GStTvVCLJTwIZAWV01UxIfHt6uUJyNAgalQKAx+N/fIYTOhOP3iucBxk+weTMJM1STozgTAbLv5L
JTUG5cCEeYqsgVeIaMN3Ymi7e0DFjc82GbbT2Ym0+hl6aWCcm5aCPD8UPP2DZQi76D6sArUKd1R/
Pfi3SWiT9ZmH/GIcWLDXLDb92NlDYiJtH6obnGgLQ5M+81afr+nL2vFr9zAcZTjv0t5nV3pBmKR5
2BH7mw+8BsE9qaw0fN3dlVaQ35zpXpc3kZslonyNmE8/pA6904Y8T4TQNu+z9gRHpyhBzw75Jumy
Z8WG1kuqMq95Ro+JeWf2jB8CYv9AhfJF/PrA1oH1soTkQrC8go7iC82GHaI5hJIn+4oc/Ifh+WW4
gxx0NbEN5NCVBev3zg4EGGhrLB6G44kUuD/0LmIsvU02RubNRVGfHaVq7HMmheeKkw3jU3TpbZp3
iehGh8LlVx4rq2zB0VnAo7NSGyspKsG4IfkIomTWIHpMp7Ei3Ga37vZESRPtvJBXaWyllPrVfEEc
iy3DWmGIMW26X87e7OnsJmivmq/9fC429NioHNu63YIl7kqcWUg89JMs5udewfi+3ey24C9VhAZS
eR2LDJvob27K7tzkdEddlBFInIsFpDWaAmZX+VkdSgY2A4ekmwR63LXSTLKc8OlmRZHF/KICGbaf
PLMIXxWJEi2z96q5AL+fnWShq4l21yLaiQhxi3JxFG+hFLiid/TmL66ioWbzli8BD6rY+T8Foh9q
Q8NtR/kBpIjDAQNR8sj1fgrK1APmZjkKawuK9kE0LEFZXEw1IEajfruXjhvJHyDO3Q9o6gygnDoa
KzG0xchv1HRgj8WWaONHzZYZdXlBTeXM614Bw5y3AUwv7dyKj2mK9iYVqpGMie2TzshcFFZHRS51
GkhD9yhv3Ifwvg1qiHipF8zFbXEoPqA6C1Sy0v+sT6y1CtqtdRQj4DoGSKf6WwuhmJjUFTiy+USG
8FDKldcrlY3QBe5xvrGobJ6UzrEqQZ1q9PScq7APUOa5YUX0lGjyAPbNC8de0Lgs1EgK6Id+prZR
yu90pKf0G1FMJ+j4O1jnYzMFD9DyZXedAmfGL91dQxFvmIcrn+qw9+RUcbu5x4WM+QB1Iz9xL7qp
Suq8lu/SkoLGMXndk+IqZNBsVmEaUQSU76NkpdwfBYIe1l13/hFVaYGwzffnKgOTkbe6UiW+2kEP
sSmGneMQl2i4+5D5W1flr/mFCT5J0SSZLarbFF2DVXjVfwK+hklGVVCe80MLWbb52n7biyu/hcU2
jHi8Km/JSprh8/76mGOeJPOBoawmz5YF6rmCMhpBUWYEouNOOgHxekB2DEI38ZE26lZ/FWSVmK6G
HRpzUDhaSkzFHDsVWUOhdLEIfus3DZZWJgzlaCbcyeQv/CVaxucJFtOUsK4cjpQsnwnIveG8G/8P
KxuLDEcxnoQlTN8dJdTkr+iTXNq07dJgw151XHSLFkFQuXXo7SdIzbMwLwDR9Gh7Ekk+qY+ur5UV
nvYunIGRSsx2I2PWd1vsffCkLFbXc3FWQnYAFmLc5GJbv5N0ykQSS0JoJ9sqDWw0Guv3WYiL19NJ
2e0HyEFZTfbgKlXLJqI5CZYJP05DkIGILRNVIvqmg9J16WJMLh6K2EGsQBzl8JBVagPmf1jRsyf1
svdof8aPpECLk3nPEMmVQAm/YNzYQaYYpyMTQXCnYE7IQf+8JTzIJVO4nQRqEY3c9ubVArYif1gr
NLaMijxT+yFA/XVoYtRa4wRB7z4S1g5gD5ly8M7mGR5kLDKcToXEgIfePRAxGM4A1fI+W/nm2Tgo
oruVDoOTq274nbc6iko3UBdSvde5pfpsboe9U01pHOaPRCIdSw0sjxB3bqTXuNlR8Tvv5NAD57yV
ST56p4yuCTHo0DZfc4opnTaIl0gZUrtlRI/3VJ+HKtK0k0o7FVdpMf6oq+3RlKSARl7Yf6esomg6
w63P9lit17LP2STVdmUG6ZEAq//Fmn/efr7QtzB8bgGKLN6ZjdB8YZtBzuQBGrjppI8v1f46uRGF
qX0MJTC+g5+jK9lr3O46iC/TT9MuPJlSYJfbJJ5WocFn9EOlKD7z60wW9mnyVyaiNNr53+st2nMV
+EqVn72C3XE3UtoMDfl9J/6U5+XTuS76A/v2xxC2b+8VYPMRBDTC/U4mHjgyM6Mj5GQhKK7ecId7
U+CoN8dYATTYgYYx1zZn9heKdyAupojo2QaWzB9jgtkxgWt7aaOgl91WBITKnvY9ZW4KmThokzA3
bQxaibP8nd45SdciuRyKIgBKZloNHYf+qYKRVV13f8DITTAu7eU01IjUBO4N7j7w3CaxKwflwGR4
qe8wGqNcrpe10/RF6wJRF1P+koz1I9vtubuJPGEn5UQroRrPePMVTaaXnrjaXBsh5SzsRuntLAtd
BGBNraPftaPvG//yrUXc5jfXw5RqOG2FjYFLvz4HQmKmdvKhGDDUtyxRt5EKJkVL30NS07D4ZhFc
2XuEJPLA3Lz5X85g5y+UdcW7Wg23rUtG6vIMeUDOoSPAVbjgtH1DCDhDgdNLpU33IGMVbsRukP4i
5D18whyCUS/hEIk6rjvyE6Nx8+sSoeFYoXFvVK6nBFGcU5PdJaGS0mNNOzPhL/q7GIV33hssVgO0
ijfX3Wubfb8r7HlvdHrxLmm2AaIMoPPstYsOqixlkalfZnmeT0LvZfkwiaX2NIBFLypeV9kDOgwA
4eA+/Uu1ZhCyGijmYXhI/hYteNlZyHTl50n1NHV1sEKawgVvphEZegjQdhnPwked+k+FI7/PLU7f
ZaiTCA+pV5esSJcQOE9x9j+of8HlbK/sv08sFxm1nwNRNmSGBdQY/U0friQcvTaaB79Tpj1aqPjT
ZC+bAsKXtPEvuomy5QxZNw/9rmIEw04FVuWM7pABPHjjOTb4BHSjIdFhfFeTIMM6nJB2YpjOj9GI
wOKaYUKySLWfxMYOvy57h0Ukv028xItVkQ/YbHRNF0VuBZ+2Qobhr5NpOdYvYTnx2A/L7k+Dr0pM
UrTgr860ATzcI1cWLBVB8KFLQUbP8HWe/50EpRzIQUcwhVLFEPF6aF65FNVjUA+Wa61lPD8oFX2Q
cxH0WpnLhEHkhSf2BOTYiH6S8R+906115uWtudFVeEpVGAysJZ0EE+QRs5Wgrg+HklBdOk/LYKRK
9NeAU46/aUnLkM4n2edAQm2K0Csta8J0RWJV6H3Iw1IwpiM1a/T4vcdlAE7noqvIJ9XKhzltO4cS
UtAvF7XLjVJW2cXs0K3Abzx9T4JZ9Z6OtjvFmjmz94e7sPWQkcYFJFqNqPwsyDD/WQXnY0e0X+ha
tufzIlcoA8OfAe35DHgW790tx3EeOjuds3rC+ggtnfui6R7vI/4Y+LtPFPZbwG/9CFytloRIYDLo
G9ePrQSpP8/+lbe6Z2C6zqx1MXSsPJw5nNFOgyGj9xtOKZgV2zGTf/CSZJom4BIGHZxY+5cJv0Gc
ws62sdybPH4tJi/BatScBTz8O39aAQr50Z/T4Mr7tTmNp/FyjpDP2kyduHYQLPNzJ2KzcmLgAEgm
Zom42jDclnld8vktMWfAWdXIt2nlrgyt86zWilqhOyy2EkaFwRG83x33CLPaMhda8b8n3K0ab3mF
NZt4OP4lfkFLR5emlIc6QzRMWPoKHeklW11rw/YSFfvMAnlD/X5zy8eQsmyfBEUZ/3zNRoBz5sFw
PkHhWGCNf5DbpyFxB0sn8UYfGFbwIxhVTlnzPraUkW/onK7nQtLJebs/x3EkasudMejs5lAwqKaV
pQFpAD4pf0HZPx4hrO1DHATp9lGDSkW29VfliltBd622t1GMqmaxu03onzQRT64Giqe/Fgh31C0b
/c7gSjd+dWqT0nRzHD/8ekp2BhJdiiA+HUmA38qyGITH0vZt4r8bPHv1a52ZpdiFyhOAEVNukhfD
s608jwQkDTEmg7f9khAlkyIzYYHBSCypTIFKAoFf1P0h50NVO7ebqCNfwc6Uo6z9youD5wS5ht4W
nntdliGRlnvvOSNXr9pvBQCm8adTqSjgENqGD4NsGjtr0BBEahFwc4QJOfnFS4cuHQXWEQLd9A9k
EcUqiSXEK2Uj10K7oBsoEGKuob4Ur95v5SqpiEhRrSy7tmuAaJq7UVT5F3+CahQaNyqSi8mskS5d
9tFIHUrr6jdw7bW9qY66nob++LZWDo1d1tNb2/6/xPfQa3DRsR7BEY/4LhUOtGTH3zjOE8t03zUs
1IatTBly6FcTCYCQILETuOjCSReElI9zRf1hpcG//41IvXPYQcPLI/T5yxP0x2fSCJt+KMeuIvog
HgP8DiMPTdOtUxnla6DRDZPiH/pK7Gi2zNrvbrzfaYGbNiwgI+4KvZOQBV6TFqHqEE831G3Gyw1q
LiiiSZo/KUMmFtRhDQ71rtdcAnBdQrRNq267gXgaIC1342qzJz10+DIH1wyMYS0ZFoywGGedPlYU
4kSkDc2usSzs13Gwv2GbOtnx8cC5AEaXEIb4K/3Hezy2JTrqjuU7JkPobJuGnUd1d4mIBHnfyiep
Os4ZDW+ebhuQZ/O/9qDun7Ys63l7eK6nxTr9Fpm2dcr+vFNPUXYWSoraMY8c7ffX1ryIHUuB88L9
VeCEP2nNKFzN70lwSt6uzr9zdXA5Mcr0y6sdqz4SOa9oDUZdYwMlozyJeCU6tIs2VrFKMJBnXdsv
lL12ACgOUguxUsvCTT51CbVks6C+L6NreHMT/SNykD4dnOzd6qpkSLSP/ieWKd6Sf1HSN+UNHm5S
g/F3echVdD8v5DwiAq7RofrxHvL2+2gjV3ccQEvmTQFeBfTABORBlZ6yTSPDdx0M69qWuOBCLHTc
Uo/hRSbf/VMdwVxRGaljCHv7We5l3hIg//FXrMB5QlO/u48YHd2UlT0phwsU/7eat4GYACCX/pu+
Ordp1dqQP6GbtgGpxccQDjymEUQrMioRpRosCsx3qQygV4S3aHzfa3oLJeLVvfdVRfl6mxRMaA3T
NVOa57lK2PZihROLBFjaWH4+/0vq9XUd2fED59ab/AmCRomIik3UNyueRm5KijRodVdPZKc+josN
6APnraE1InIRdwjlkn0uSKoDbuxHbC+plg2cxuQKB7SaRMDhQuOvrXWW1Z6r1uzdQjcp/2sZWiVf
QKa3dZtSN8BKq/y9gx0tN5i9Wt1cCtcb/V20DUfw6UYDwMwEGOfS30SQVt2/nCprLgcUcYgoPeKR
mrd/9TpTPErdGNqlIVFYrqvh6Tsvl8YzxzAK4Y3WeG9ufOT5XBYS5aVHwVqEMubPR2gFH5qjJE+j
KChGmtt+cGcKPusckkZEIMqdMo1bzamE3uwNv1lZgQEH/mFX5Rj0qaeZ7gJXceMlGDW3++XzM76G
d6KWMPdhpD13mslqMFjpl/fDybO1NILyeLdR9CaMUsQxwICLHnbvD3Mb1VHshBuSAV6mq3eA6pzj
KdhuFatIxPX21EsjwLw6qJQBy1CDMQXUE4mewMYQOu5B/P21iCI6xENgEi1DUr76DxaPFDPCwLon
mFmbyJPEA/WxVYc/Q7m1B9mBEKKP8uf+WRWSCEyhQ6+WRGcyXRsBao6y4iYX8wZNwkiPmdCUv5xu
c48LrgW8cefGq6Q6IuA3y/9MQDszHzexcUAOyYvfjtMu6fLzP5lcbfov8J5bMER/owJFt+cF2Kvj
fdjZ/vY8snMzngrrSCRJMQutWnp+cVZ/xeAbYeYDw9C6u5ZexmM9rjPOlelCFy6uOvLQccWHoi2B
R6QZo5EjG+ViMoXEmdolSlN6wJxToI0xvwNpTrJd8u95MEc9gnO5JydqKGHe9TZZcTS+HeaOyNMa
kU4iffNKjnLE26J75s00FduFOITbbIr2sUYmzdQJKpFZIZ90ZYMWsChI2F7tzArlseWbgr7W5t6k
Ac9NoknOsVq1KeTIZ85BcSUtHg5mrDpX6DICwNrzcDdntLQp32BqqkRagoUGl2t0I/h7mM2E9tKp
kowJO2pyLqbd1vhn0c3kxLVeIFop0PqpLAnmUjIKXesKqISKG8bMx7HR302bB3yWPWaDxXQJ2kha
2JgxBK+x87fAE0NgiSoxVqAnMVygmVhfvMIk34bz9F2jHz/kZlkpqanTjvmrD/q9+a0NZxivORa4
DsVjIRFknCzNtvWbi2GPxN3Hg7KK0recWHb8VjwKCboBLeHcNFObx8hm9uLjc6ZXW6lumfONfUm3
Cw5LXABYOmoWShF+7Yof7VMRyegzl1Emjx+6OBXmmBtnah3EjsbtyqBxViQiAvDBhB+q5OKKDnnw
hTms7ggoAsSWXOx/saEr2PNCJ4U3RhmjRy3U25IYuXegbq/DDGxJn1uL9e60CRZ9r5hmPjQvWWkK
gk9l5KEXCcbwXP8iVwdtAwR8C56JOnGHDN4clPCKTvgEirHZvK52/wo6loqgi/VDC1dlSpFv7Gx4
KQrw0O4VlhkZqjnvu1jFUTRm693Ku5ya4h1t1SjTCA0v7gIECJq4IDoZS/cBLc65Xc3nydAx/fEP
Xb5CoEXkzAS1jW8YR0vG7+CbvFa2ovDs8lSGyRBFtv8GzQCKp5H3fu8HcqZ8nvsAq00/CjJBZCET
DkVkWn2hdRUgC3SZYAQznv4lKj/At/2TvJ0h1hbLBLVBmGJw9q0oO5IUPCLYLxHM+brzMXRiDgMU
K3cbN/PXNJe/OTZ7Mj8GGX5BBlKrHPKMd12C1aM46v4KBTZiEBnPD8gcl0iISC3ocHtQ1vSm9YJ/
PTmcGshRqYp5UR+16lxe5Xw0YIuCggmmygEzRWnexM8eu0GSHTqnHRZV4BxBVtGFs3N+/df+RrK7
4gDltkzWhllzl0wY5vgq34kU0nWE+WqYZQUwdO35Ih9FQGTlh9JGObjgnaf2Q4jiKFNu67YDzLgU
azMEVepbpTOcwC1MYbF1b1Q1/YQjpFoP34AAnV4usN8gx4hcIhBnx4dua7KiJn5waKsSqNhGn4ag
hekpsouds3NAP4We3N2rseNjg63yAUgrRrT7wvbsC5v40aUZqZTYTiye7YpB5PE6jXjgn9OHbktM
pksFuM2kVahmpcBlFs/WbEDFpvFiLY6ryEELmdWAB7haTCw07HNe6qmxdkms5rPJ4P43cLO89TPc
BuSu7bcT7P2L+ek5k57E2p7XGTq45c6V5uRWjHBE3VFVWI1pbFgHOCoQUJ/N2O2cDN/Zb3WAVe7i
XD9V7Tg6v51/wnr3h4/+FMCAs0fyMb8rcnswUehWSWz30uM8YKa+FnghGvjW0kD1N03Ne/34bGQx
rumcTKd8+Gl8qhdeX4oCAdrpsm0FUerkb2MOYmx+iH1JCUOCGMPea9nI9kWHwWtc1TQi8VKCMiOf
YkVoCARKlfe5mYNhlVlzTTM7Fll3bHcfjG25hXoV/eYRd5d64JPXUwDHaAJttpnOBycybVdVdYY1
gnHzNFwABye2F3NhVFaEgQU9VySiT99KqSyGgGK8ia2syOIWs/lNkLLaz5v9e8rKJdvdiFmx7DNm
Utqi6c4D+RpycjItiwb3mL6GgiU2cUbhEjPx39zMlq4uDQOUW5s821uO3Ghx2HgFwhOnP76ZARsZ
A2ILPw9SAyWNCK2QMGqVFyMvxaSlH8NvEfbuqGyLZ5x40PJQKqVEv+MeYDhabk5O3nm0rpU8qJ5v
gxO1alxt5tTsoiPHwLvtJEQjg26rkZfEZ7eqzluSw+60qEu0SYjTZHBkbp2Un5tP+MSaX7X1589c
KMRxuLeuI2Ju/yWicgV+NNhMaGdrIzfbpLtnpY0Ex4m7zHZu4QXEAkqNkbPfm5reYEK7aAthgxkO
m/LM8Sxr+LvqGJrsEtcS8eeiS7dkBH+RO7LnNEFKa7HbKNW3qbHJqGSmzubDuSfHR6LMPPdyFCL6
YKd/y4u/5Hppw2cQaQTBTSY6S2m9vthpAVLQgZ7TrLsd/3kLNXzR/GHbTyQ0AvI0T/8DRAbwjg9r
fGV0P4a6x77hX5YTnY6RuTa8X17H4nFTWSIlLWDHiCBnbjXYDS8FHKUMRktVtpbnGClw7OmFT5ou
Rl0MtfMUPPeJ48pmW/1yJAGCCO9BviHHi4j1EYV6yDiSTMnGuTLTLeCpnSrd/4KSesi5HMwF75zF
v3cuEJkxYhmeEnLtkrL+T1etBJ9r99slPUMofPXjH01sNCZ3ovUF9vceZjyDRQqJujkBN2aVksQm
2TXhvQ3Azq86geoWR8everp8fFyEF1u/W/xeN95vDIMyrnEk2w1XfWdX5D1NHwi4bbKzQkqp4x32
ygDNMYPudWYL3kmqPrLoSTCYqZBFgsnBS1TuZUoBgQB2HmHD6TSAP7V13mNQltm5MW7dqjVbUhxI
9WhDraZrr4TKHS0iNe4CalqowkPg50s0C4ONjC/2eFP4CnVjYrDvGaBvdWiOhwfDsCLk7FcriOTF
6CJvWZF9hJ9bQlFTqTA5VoMclmN7kpAElNcfAVZbn4Rhl41Ej4XanuvgaFrR/u3XG4M2bTx0zODW
YOuX7NkEisVlBxZcG3vCb1HLSePiLrWaw1EQSparMvGZcbFFGknEp1xL4xdCgFYj8ASky1b3IL53
Hj5H94aC6e2pD90shtQy8v6m1g7MZYc/YI42cdxnNxbaumaE4gI4k+I6EUI4s4tdXZYBLVEzMQN4
9OJEwfWBVmgKTxnv/KsNe/3U15IQbE20MvR8zEsLqHcgU6Z/xPk5rNWgZmFRxKsiyzBCeCNRBv1b
mMIM7Oe6k0GiKYPoLfPY48SD0Yz8KN5FLht1NHdyelrJttuzv/pww/C4fHHnOXWQl16ebNw0Ea3/
spdV0700LVkmmsgFMnUfpsQPyomggG3i8aMsEuMtpPK90Xopw8Prt9oTX/AI1gE3vDwH5MquX4vx
LoihLI/MjFZDHdIa3bvq/AEd5nVtzo6f00kNq+ETPVgeZZ38gM2savNer3/aBasVTGfSuchZ0G2n
SqNLPFU1I22nMfOLtBCDzM+bQ9z83EShgpirip/+uRTT1T6ndlapCbC7VYxI2Rb3HPtxlriCtJC8
x17xdCZ7j+gFqwJy+HfPh4Oab0N3gWfJ4o5XVQZclbkb1oiwlWyFHINC5xOOtlDTdK1WUUXJhE+Z
yszbLNb8N7eJfeRCr7nCkpfNbG7gYyq17I26YTN7AyoU0st6wWDPI533LuF9W+pTfDEpTGR/JUFG
rSlhhmY8re2Sh9oRbhFyTV02V/kurRLq2n5OBbH0NGwzbOPXmeWF2C0esOqEUg2l8QfAFKY403w3
mY/b8v4y+MAHrqTuBGab9G4zR6CbmJbBwS/m7Zf9n9t389/TafXEpvjg9XXcFI70nC0jB9dxJhEp
bTzP7qG07ZwSqM7HLNh74Tmi9YWi0TepN4MyGhHrYKWmYoAKbVLlP8rK3RSfiScT/ezCNyuTVtbD
3EDO1z0qx4BQoiXSs6g7GcH3LEYz5LEQzWtFTotR9LqidL+tznPrfiK+kAkyFHvXRcZCFq0iEFEz
ElyhQh7sDgVMkvsq2dwoG2YKUCyNjJXUdTqcQaa8Zg2PRtjcZZeuWBhhUIuQyzx+zAzFTAXHQibM
+goNeI7DGaSmh1OdWEYwikI4cVNkX8zk6tacfrxm+BnKj01YYQPDwhKc8dU0Eajv75CUzEa/F3os
h+WxW5jz/WdlTPzhBfpqOjLEdm6BuYWkFTiHz9h7x7mUbu/toq9ug4/aPg6cULPH28XdFDZWPNLy
9QtxjelGmjZVxab+va6/b88pOefNuVvq/GBbHxXTcQxHBEZ+tTg1JsTfejM5PgL1kTWnY829+ao0
1jd7GXNVbtN/arA+OsDd+TX5QZeLIukFam9fUs/QdIKEfhBP7UA8ylysoJ2ONbWHFW4c65vIwQlR
4sMqXbeMG9mdCuV5hACigmHBfaV3UxcbEkQ7Z7OHK6T7JN1/LQNydQavu+prwOIvYy75fEjFtfXg
Wd+lBfm8Og3RsVHLLwyJCAN1Gs911bBttpC5Uy8vyYKUkpWvmYa71sc71YcpObGlOQeZrMmQ9Ym2
cf1y3jDXuwbxidb+yV4rGshAjWyiF26AyBJDFTWJ3BWXH8QHWJA7wkzptE7l6umzCGX654fupyXg
LwQlod0jgGu4aF6x+cCzIWkDrrbvNfFkNRQSB0RqMvQsWjyY6V4W03m1RHLa28ycrJ63mqbqM3cK
MDZH7X0g6D3zvkOxONW2hdj0Xyqkozqng9g/GqgGq/p8ItJaEIwGDrIyYYj6dk2MoEit5aQLbNLL
G46OYQtAMRrKeh+6WIF89dk8FVfg015FN32jN5TZrPhq0LOC3NGyiqipJ2YmwkrX10uFMmzOvHcy
VfhmL4J07iDKboUU82eEvDiyMNJhsO7zvOm5iLaERI204oNWxSub45w9pFiujrhajbEg58UzuQl0
KPeouRgg41h8jp3fP/X1TXCdnB2ZVtwAzuklA3z4m/7aPdbgM9Oyb6B/2gxnABuyFDjACwJ72lVL
Cw4UHiE4E8Lki0/Ndr8Gz84+a0Wr99dHTQhutgGaMsk4h3ZME5ZH+YgGsl+x8ozSbylq0B07zNpr
7vv5otwDAN6rYigkerm4AdfAEgUt3JKMVGwfw8gD/X8tFphPYb1UrEU0eFi6n+NNS9utpGf7R9OD
fRArsKGawg2q7FycXR0S/63FGVd59bfYwJTxTe40N9IZVeYmNL2J9ljgzaQ6Wq/Ih6vuPphjJPSQ
gn6oteEQLPxRY6By9mbOqaoeMJ+49a6wAtv18QCxewJguK/mfIym2Dht9FiEX9pl51TuXLtcJZjX
uFJ49tVffUhZW+yuwdsdgVMk/pAUwrjhpUcP7D+3ZQiUgDr6FdGGsMz9esNzpRyUmlB6qdoV1tNK
NUJ79JPnUZzQ1hi8s21qLke6QXFGxCHWBdIhFuNIaL5T+L6W4TuEXCWh80T4UBkBtPTfxfCNlC0Q
NTvQV3lZ/6da2EqJYBVSGdewStj1H39h6f+Cbc1X8c6d6U84Iy4WoWTbb51bCYQyjlaVXCremrBw
hPfv0r4KdxHFo9N1wmcwecdx84ZbVvoU64eGOckEAbXwdMRc6kjPzQ3gGWliGVVn+0YEQONB5rCk
uyjzT0tU+rRkr7E2nUXSs+wLkBF+VtZ5rjsdu3Ys7vsqI9wzhiU9o3G5j/RhJ0QoYSaRPtTHC2ST
kzvl3E+6c5fCiE7bYMURjWk/D998ldNtGf0ybsaCP9PeOPgr0GG7IQ0B044g/Cgj99FMFHEJoPcE
RsT2Pld4COblafJY0cyS+FGd1L5hmdAzqYqbw+ug4DwTuHjZ46/unSAhdR3TvNNPeEuKtDpG0Fju
tFcEBHjJWgHu+kw4WWrVjLzEvfE4XEXSu6ADopYHdUS1r03Ikw+oZU7K8MkHtz6yvid6A3I42uhN
X9T0G2LAccL5DvpX/NPQ0SCwcrEgMmf8Pu80kxRMXl8flbJI5GsREAKzEly+0DT7b94Ghpukwp73
9huAw29pr8lM2O8R+NJ9Li4xFj9b07J2Bvpltyg6TjFQDFy4JeSku67PSZEAPCKAzyrDdb0nCoDT
BwUyNJ/A0oExgD7ViyQqnLMVlfVbahzWzi8EMZB3hr0Bi9Dw9hxJm3MObb0/lepu/WJV9PflkGk8
CMzzFPoU3a8CXceNl6B10Abv9s6QjudtBDsLJjH/N7KFIcILUDRisNaikUZJTgZwe9VuecWX6/5z
/krhFUrM+1l5VTUAonkSCuaj6WwItYiGwUEpvYQpKxGy8isNaQG4nZKomzlqVY9Xa1eMlCk6NuQ9
u7eAdOOCmjW2nIVyyMAZ+Cdc/V4Dd9FuOElXXbOGVsXMraWLxFSh8ZpmX5yiPlEvYJk43WRic4b9
dIIOTS1YFXxILxovIDYUH2I/Au5QC3kGVKjlKlXgUj6GeFeMRWYmrINR/+nYEMcVQK0AMcZ5gGsJ
7ft8cQtztpH6nKVmqd8JVbAjnPVa+zLdMX2DPPg+vUKCHqmb9uVDAYvs9hgjctHeFzp0UkOvcQqn
EtbvuHZKTUulvWbdeE3cqdhEkNAtNRtXyZQPpVU+BYFhlfO83FDAwW+PfruFvDcOkK0inlpMIc8F
N/nyQ9cD1FumKaHzayFdSsiu//U+jeXQ6ou4HXWlreYrvqD8kj73LY8fGbsy7vozoMrd3FfE+JFe
3BXNTZ2hBc/0T5yIMX4NA/8gyBKZS4NJfjozb0cABE748k3wnsa93pHBLLrhlaw4XwcEo9ZDyic7
beFMqRSciZIiUvUjK0vYy87MNtNQJALK+pCd43qpdBPjSjxbuW6WWJ3o5LWAcJmZqqFNWMeV5Il+
m9GsTjmEX0D60GsSWfTUyse8xkHJ8cNS8KUfPntXXgkyUeYEHsk6onLbvvIMjwh6HroznEBwrXdb
YejSKRDiJeNktB1Qnps2CHLnNZrjw3h/Zuf0m92xCFNIw7WypPnruaprwBoXPB6KEYhTEQOaUmoO
GqiDAlMO+NbVV/xEanv3dGWM49Cwd74hWFJSIcoiAlQnUNRi+FAHzlvNepxgTOyxcfu5dUfGS6tw
QKGp5FMcZpsGT7ObuxHhZV59Pe2HfrtKsa73jzZbTmZ3p3QWTKeQYC8BP8tIlKP+t7wyyCVxy0Vh
ioed+8wBKV5zIXu4HgRQnJOnPrSQULfHP/hu4LYpVGZgzheY4z5d5j1J+8eXpMCdmSVbhiAjOTGv
ZOTjdKWWiHjtQGajkBrniJDvMdtDmzfo3wMhUajdpMU1cBC5QHGQ3D+lqI/HadvQYwgf3DBq7P5r
4P0ubLBjLNCuU5oWNSrrecJCovPmsVS64k6yyU946FoKHMVvtlcBoeX/uBa0mmMFM5ZivGTILBN4
xt0RCR1WNNN7OB8rrgIua6mT+cPDr+dm+q+pGCSaGKOyHxYDeJQWlYFiy8R/DoVZ0GdzexRYwYj4
EUx4nZYmP0lmCx6wfsuJ1mjZsqg9ilDAX28gIVkYxV+ljihNK/tXmVhUwP8PREEejAgL8B48Hohg
kVw1bpf7RfVTCqKOFSPujPH+f0+KIR/s1J4DKpL0kl3RZ+n4GJdpQZT0wInn9P+iwqkL32XXJxsJ
BALTLqfdDW3qfTziEaE0xi+6stTPOuk/PBS7BjimdBFO1uCKYVM4a7u1Z+r0me+tsC5gm6iwnsJZ
CEV7dpfa8B4RSjUnKWCNatZQLov6/I7igENPh5XUzBgCqR95emQp4s7tKYK5ZgMSM9LvUeevdC9a
o5OAW+iRhuuC83JC/oIpBbczM2cmGaEK5ymzlfprAfwgz4kiSLcjrvCCCHndqNrjOYtcYgEUN41x
IJjMwG6AvsM6xELKbKIkoeyZpWhqiY+KRHGo+LI1Yj4nGwiVF3xYxqAPwfHPbi6ZoEjYftDRYGDp
hmsaqpX1FkJdPJFS9u8o9zzg4kCCJFYgV2VpyfsNPR6wS/tsMEQXpwcQhhHZOMH2BxQi17Lhu4MR
sXq/XAn6jr7Bvdj/wuxR8uwH3t9b2ZhmSfRL8zrDVwLBSTo1iuqDTE4ePgCUKm/VByE08RVkYVZ1
deU87MGfsB5/CnpMFi8UQ4nIqJaz5+D0JgrwZbeOBvQGzt/UKLUZ1pBTrnmB1S+ydzYg7P4URpEp
4DJ1Mxn16nklpOjOfLfU4gvShjDgcU8ny4iZ7rr54ucoYs30HcyX0t9zfq2Zqq4pgJodMD8QR8uc
v6wb5j4tJavNteogAy7XC3mhOyeOvDmxLThPbnuM+VWCERtbImUFG4hw907JDzox7gmhv/3rg76b
v8MLQBjz4tm6yYiD7SmNeBNDEJ+zdPLY/TToPAefwqY3yaKbZtO4deZ9HZ2JiHJvqkaTAW9Z2ZUD
RB1FtEsJJJ9TPIXl6j5073f45EEv7eSoFWZnCcX9xO2WOPD55mC7FEdEOIHr/XlGzXqfehBXA43z
GrqSMu7uC95IdADXSNOdNVYK5hoC3Xgh00oOYBa9M+sNqy+ljuPNJYAAtNZAYZJH75lW6SsZP1mE
2EuF82TLGLX/u8gQfQvZ4LaMfrL5HEL+SL2t4lVWa70TUKZtbc1AWabiLC8XfpDFh62KSzFbQbMZ
/P3aW6uz2h+enz3oiWZj0AC16UrIUP9ViiEuluwEqnAs/w0WDcSXVMHqwyJlBxyAMXMRwCh0cL7W
lzkjpSaN4tyXN/TqeFcLnmwteeCDlc8PK377BZJk/grm8k2KWwGA6NhFPzJ2L8YVWxLVHsCxwAd/
7WhJZXADK9vDeMuwVL06ARFsIiIIshf+TD8HaEWHAhxh+ht0E2U/XUzPEQdrrdFTHFABRUyHGVhM
ajaftTcPMOWk1fiUyXZcIUyk96+rw3FhbCFFuyhUyz03BOqLP+gcyvCluh1U95FSBLRxjaRK1LlT
v0jtkFRBM7PlIGeTFMDoj1NEUBxjQJ49tkMSXV5foUm5aCtaUA8yYA1LfsLDjRldtiXvRoG5blkQ
JeVH2bxiZKp/02BSL41qlSOGCCe2pTGXOpxpBTXxqhpsShrJ9YdZwRCkWHH3Z15L4g0nvau4d0EN
gf6aW4CNacgC+oZG1+2hjb6W8krJI9OzTTqdYFDBfhCUeJxr8qSWpHB3KrAEjVNj8G7ingyvTb3Y
iKM8QLoK3Necfr+eY2x7DO4U57cmhD8dD5WrD1I9vy0zPGSaPcZKNdyi3BHzZ8ytOGVTt3ZC3FKB
sPX2ITs5qoxoskHCuYXeyEEtyMhS5TSdl40n0DYAtenkfOKVvqAd1LItSQncqr0O+kUk80hSEEYH
qtlciSRRSQeydr0TXivF2zGB44Uc/cBC0UdRvKnr3NPmcetgMN/BArsPBD8ugZagWrNJDW4KQcxZ
u2D4fxA3FkoP9hzI8jbb1xAqYCtqztuUHxgD2GOxrYlvq4xvXWGXYCI0s3F2YgWYNP4hvA9GdQCi
kIrxDXBKYe2VZSZRi7BKcl8e0qbLQgUSk5ZF38VrraLdQYxViyiptR+nDs3fKI4Acq4dl099rsAf
EqpsAocEehwZYg/MaunqQMj2U4AS/eN/q150SLBe9KiLiF+dygN6aGgWHbYFZM4+lvMbo3AyXEtr
fy8qxyGKp8XQMQGFvf15T1RMOBKWIsR+cc2myVTewiUPtMVk+al7jZzWLzEa3ov8FspcME+fKxxl
7OXV4eKmX0dL3h8jiT02cgQKqLapLt8ubnKrhBf3+jjdD8mVNIYBcF6hkjgdorc/bdcDKPWiWBMZ
0MpalQj9ezn/s+Qf0vaWeWNvfGNgKEWwOgFHaQO2ScRQ1d515VMr0FKUmu1wanW/YIEKBxZxSFgT
Oqhxi6X0Zz9YHAhqdWJ+IY9gBtd9B7wcr0UEPp2oPs6oF0bUj+VDc/bb906JlQlz7QNDsrrRz/3V
qFuLbFgG/yOY4/E7FhMuILNkW72+BxTTvfkBklS7oaDFLi+pbgiez2CQoEcD8CL0a9t3tlM69q5L
mphMutN9kMzDSmZ4c3gBnvjdNFOlwPuw4V5jU2v9lIVdxF2lJcoozv1zW1f50/KuJigwdLv1iLMX
+RpSn/yTDRrUr7Cp6nCDwqvjNMFDxd3KO1VQoBqElI291omO7cvPT0vNeTuUqVpQeHk81YkzcuYD
HhMw8loUB+YCRMpesc2EuzrG46FliAS53S8q4fjfLsKVu0PRm98OSzX8olm+KogEtjV2OUGhN2Ly
DggUUv+U8tD3I5m3DHKEFEuTyl8p0uCIN+NThCwmpfAH/KeIFVhIOl9lgJJL7yQn6WdpuljSSyPE
dnb8Oo3XU4TPLCH6f+px9j5KMYpVQbOCZh3YZMvI5To5n+HGRPniOV1AReZYjfZDZrXYRanCAAYH
pJT49nU5WpRbGqo7K+vV6CJrsHhkJLJxn/ckajW9DkFz/4pY2G1NFjxPs0KhzkhCtn7TqlT/SFCY
CmWLHSPufub5yK8hl8KVjxNRrp60mDgmOxz0esObdI0qNAZuKYUtZRVxuaeJYPnOHZ0sAZt51jex
9oFR9RcaBt93eMF6XK/99iIMr1QD7O63LNDSIG7Wd2hHAPhnQ9IFQurjKSigseDSQmUKCFue89F/
R+oXXJsLwhLzTzXAsNiILBOgsjgi1k1zhJETf+O8cbT0ajq/1Cs/SDkX5etnEFv2GqhUiWBB5+Sl
kwIlDLQ8h7gCuPl/KhiqzS/Y2xCJvhRu7U3ORvgbR1aiRahcu1hpLOGwnss5p/AoH9C75/s3sNy8
xH8gfJB7IOpqjeEzoUxb/vjmWACUrliW5Ww2zwj0GzsA5+XpPGvnF9XOJ9/jqwxMIf5wU12fEnxI
kLadhByDUBIWS9bp32O5tEQoqUrVQ6TTau3C/98UcsQtqv7456JCLxhLTd/PiPV6DWs3q2lk7ndu
YD0YLFXmOs4qkLlTaVq+MGE6tt9pmEHENDNuHOxz2ULiogm57iVUN4dW1wRRSxhoQrkXlU2zGne3
BqDuZq9b4Fz2ytmYl+WE7lJITyq7Ptcp4BwN0kcpRK7DuITHVGohWmpgIq/psnp0GmffNCGCtSiH
SoKCSQzbjZjSu11vl3zVEuy0V7v44Wx6abzW8HO/CGRtmcOmVI1LPOnp7HO3uDuoGQIRxdajin3m
xcvIMeBFx+Wsh+/3S1T3jt41NuuiGKCSq4ik8aBxBiI09xqET8vKoIX/ehrezOlM5qoowihj1xv9
Ar2BxFNS0NOIk2rb78J5LtVOz4Wwtp8CYak6PKisZ10nS2STuo6QwAzuwnq4z0eUjdAfQCmCzm5R
Wi14w8tAsFzvnE3uTIGiq58VxQjshaaHKZ92DUlMXZ/eIyHdD0fffHj4UB/FtecTw0djiolnToDk
z2iyrWlt9YdSpZi9o6XAVJDTOpwZ6RBPNZZJyKVshzDhkLUGG+NvrcCBXSwUuh195ABSBapc18c2
rUPDFvXAXMDy73JwGeK7csUxeOb9p+mBz/7/MEkmzQD+gM59nmJkjnQzoO3eF869N50ZCmJpdKAh
vZgNAFdnn9QkIN/IjAUZfVNAXosRxEu5nZhvi8AQQ3KjJ9FsQzOzEgELB0wVgPUS1nMf7gLQ7N0m
4nwPr95ciOUJ8c+R609oQzj3WoexK6CUjhrmO3BKgTexoBojJx2Nkcb/n7CPWXrYOOKb2skFrX2O
5e7Y4CDmSDwPu+p0KIXWpVeeYTv7dpXX0oBv5lRguNN+plnndR9MdIw20sW1aBS1dOBFxiW2+djC
z8Hha9I1i9bsptQdRhP9uzkqRe7iQdNSIe5voPwr8N5w7b1xGPLyRIIy+VIpNzM6xIChbYp5V4wf
3WR3RZjoIrqlCCqqpPcHtipay2hNFMsrNCwV5ueDaHtz0JUa52lEavZAhslca/Dgov4uNb9cjK9S
4oVKy6HvIsJzFIsOD5HShywQ2qdjZsEZhatwYf8WlJWLHkLQ9ijJ8PZurawrrxjyFekON3AM6OHN
GZUyV+jd/iJS7IO6hklAcNHjc4tGebfymtvAFH1u6DfLzSpJXUZf3lClV1oIAkrV/LHI/Su2+Mdr
4lL+wDHGJX7VqeAfyHWHjxUc6Q6Jalow8j1fmRzD9otH2TOCVScqGRV8mX8KhnNK1s9ANdAvPp/4
Jl22CTUyc6mMxkz7zvscJzQ+kQr86g/hcdlyk7jpBuvQbngVMtNj6K0SGD6Wjx23sP795ZU5ezS/
pKJmA/7m9ttVED+6sDT1mfsqvT9oBvAJulpHrUZKi/BZklAf+wRKSX81y6h+66+Oi9Ycztp+2EwQ
PJdbwSumDTMlbmto+wCWcsVBhlWFuzHXfohYKLfemaFmyignywvNmtsY4ZkrjxOBeuwU112j/rP+
7zyLuqlqZsORH/NnWpA6OQ6EKkax9dnR4H4SHxYw35OmE+ogzLcDyN6LPG+LlappKBGJeWCQuwR5
9edzlnTGNxnhzj1K9uKNAi98TsTU/OSyarG0qgonWCTVO8DfpsqZHERmbnhB4jpQOUIUxQ1E8LT6
2ipvCpWWJKP5s36YLu2UFq4zqCLwDrvUxWLg9vtHWcI7SwrA5XpWExYGK8x6jCdjGUbQy7TOsf5O
zKZcLFFtgSHazvnDRh/L4qwhAtzk8JSuopVk+XnkjAQE3e+yTapkW2pkN7Byvuk9DRb+VFvQrETt
MZ7IUB16sNFFrAD/mKPI1lt9GeMqbo5qMvSwT0V3GeY05kggjbBDGM7xIWqhPLhqEGzWByFnN31k
qot48nC6Hsw31jkXzDeY668Wco79KsyBiksYRijBriyOimMVOttdKO+h2qCrBfRM7o5aArS+Jf3f
VEeJ6ADmZlbglbrkCAYXmL5lWY+ovHHS/X9M1drKDGLTq3QUESDL5V4ySBszDF1MbTPXWkkL7TgO
miKTO6U6eMI/vER8FkMenNpeymNsaSz199LeMNPyvYFKN80hCnB7V/S2FpWD/AL8Vld7T+GMWyS8
pEbusVTVjknZKO5oiuQXu5zl4uks8hZy70iBTUyf1PZzRGEsbllMjzhT+fm6K7fx+It1mNbJdAV3
qDC0g/XNtQwzpu3QzMUqa5H8gba4E657kNond5Tgne+BsZe9JZX0I+Ogqep0erAFKa3bMJxAAZau
aXmbjfaaK9Oyvjwz9knequtDbh0BUP6ldueNZ/AYcm+LbZ4yYH/o3jHV0efUm+sX/1AlwTxNUlu6
h/4OsthAW8iL4Q1Qj8CxW8PTbpn9oxrQKVrI1LL5Io3/mfZSv96hR/bCRhMVQpq2D2vWFJtegjEJ
vJd05GTa9fjn1vCVnLVcvfKha8WwtcB1hPBUBEWhlkK2g3pCUXLkrEMPftsNPIAXp/OT7sPO9C7k
dNo1d/G5sUBXupeoovudVqkmHvAu6orzfBhdXR/bj32u/UIbk2qSxjU4MUQbWevzqSSmDROp4qLH
QSYfrkKAnVBk/LANIj8z9BS5x2jXBNNfBk3HpPHMASzFw5tVCQOU/I+nrEj5kqD+67TKGDw7BwbZ
MUR/wBusIDEYW1Uw0n6fxunIvdNhcKPwx932g5UP2G2oi5MTWsO5f3yOWhghgZNwlZnizsqpD8rc
B6oJYIaIUDZJX+Oz/XmBGaURPNuf7mv00PNQouZh6WjTt4dnG1S3T7nJAEamzpBUcBw+qM0+13tz
POJcmTPU5KuSWqFqx74bP6kJzHnl9UYcZ/tNsG8EhZtNjrwiWC+8XcyMMvbvAQIUItk98J36Mz9n
Ot6YRSKIitCc9HL2jm8l5lM9eJ1Hx82KdDwixKlWzCBHMrIUJSECNE6pV6sXZMSrmGKBPQ+ae+CI
At9ZXqWV3E1n3r4tEOgdMtSaLD9FlUZo54LozvUnjs3Go89RedHGxeN7eP5mcf4LXNyI4CiwmPVq
WvOfGhX+dbElJDeGPKFe4DGnxFIs+nZuitYzZQN1bm14PiEDi9izn3O7yTn7mmshvoyva0p9Njnr
nOgu7gcPZgxtCixYXKLaoiRAa6fqIGehCjmfCUr0o7F4d/k8TOyHLwkAoEqPZK94ROXjzUqyazdX
1/lBWI6Z42wBJdNIRT9P9LfGQh22DkNb8qzDjuXyx0XxYzfUAlOxcTCdBetCloGHnsMk8AfxtxXr
iwrIbjrk9DzF206kSwKBaOH5FHWbRZVZ7+Nw6x0SAxc3Tsk9dD0WpKrQPDJawnNDDZVRnmhc93Om
EKKLKhjzyBh3mlmElaZnx6ZmovUJlVkpb0Ls7DINQrv3Q+VgL/Ov6b0m5h11aOF/Yx9VGR6un9RL
wfk0vjzyo+6KcqAqhgxN9I9oquwuTgCwaXytagr/wOvx+VlU0K3+R0RLYdIE07BwVF0s6au3eEH9
MuGUMWFK2Db2OwNf5oA8S4T5UVT3RJNnACCirzyZDpHj8WbXrXq+h0VZ7h3C33KpMNGCFzSSPeNQ
IdEwXWR3WSo1tGSe7MRyurs86RDailcGEEf9pbqXW0cTMP1Kl4PbLX0/kRtYoH3d92DJFsITAAs5
QXG3GW2QLphj2GNddd2zXZ+DeC54N0tHROFAmssX05+ta9ys2Jvf1L7DZht3qxsxxpPR29dV5O1w
934ZbO6Ed+u9Sv3KPYJWsnf3hW2oUu67B2T4S32qWBA+n+MDriRKawfwXq1Ae9UWV6UAt3AMYbZZ
LNK/DfbsT6deo3VPsGsXpcZuABUtOnt7FMme6pFTfb4ZGPZDguGSDvbSlmt1Q+rV4oV2g3ZdWPZs
pV9Z+y1Am10ng7QtrkoZsfgtTvo7HJFgbswqXUznqKiGkD73Wp4LA6mr3TMOHYwIF0ddIr/JJ1CD
9MAEmke8dpUz+xI1QT1pkQF/Eb8T5oB/nFKKrED8hmICUCQuUKMPkKfgEMJ8nIyGqgCBzPB06iTH
VjUUAwdNwHNEljnUzSOzLWL20v2TjQNwuTMX9sYXfacA5C4X8N74h6MOg1dG1NZwTn+lbXE3/2Up
XYamCyVymNbuxrK2AqkeWeC/fNm9oQha0MhRc365jxWxZi5XMBCBIb+OacZSWocIhMkmBU4dchu1
N3FqVg9JcYEpNY9KipjiRLNvad0w0x4VLHWgfjSGhA7Dd2yU/RHyXUTP+v8PuWuSkbDSeXPiY5iO
B+Ju7p+WVnIIzI2/jRdlS0qa3/pzuDLs6D5KXGVsfZTg1XWJOI0n/rrMVH/+7Z9t6FFXIfGFOW3b
vKv7b5s2PovEp48lIL8ZGHWwqhVBzH1bluXdYN7vTZ8hbI1HvLgHH8tcZ3dHfwUjrNmO4NtZ3jba
AwynPNDgbcdNATow1KYbl/HQ03A0hwMFILIO0hZoGISEXIJPfqq3evFRe5kkwkSyKOt5XVhYr2ej
4lmngFyPsV8oxPBa2b3BIQQLc4OIfwy1p3OBk0z7HtkGBM0ui4uP7pneOmtaC43ZvZZuwq9pFd//
X+9qDz5f/J23c0gKtaota9gOwfFLun6wljhJT/2AAQRHZBc+0XJ8cfgsgHPGHsD+dwghBcafVes4
PRMJq2pIaFBwm1NXWBKeOd8Q4rpAPD4fTX8KuqMxqz6BgE5uIqnLR5AIqAoOSEyBK7o29v+9Ge2x
zOQhO+qFS/mGzZOmH64jLgSVlUW1QgTW+zXvpXGdrVNgF0dnLyinQXXEe6oXi8kMLxViDOTsWiIX
i5A+VVhl7IUg4YTdwR++9YR9dTMeQs5dnVlwuMJQ92H5avOfP/ADI2R1M9tcIdJKZ9/u+c0y/IF0
Wi1Sy6OC1tYzFDcHweufi3+teDoh9fIrDQdvzNW8WVrSWFhNMin7p7yVae3AJuzQV/fEw0EFTbo4
jxe6CbZEDkMtl0GcsWq4hzKqHASShBV8A1c77L8pyN0yJ5yV6/nnssvfPg1kbz5j5lXa/ODPINor
XGcZj71AHAd85TfRTjsdDlRn+xC17ijtu3LdghkSfI4kT5N/W2SySPp0E4v2tO0F8t0OddCRCd1M
QYVwuxOUOfIh75FavL93ku7/mMI4gH/wxRncIKdC6bbPOqSwv22HNhoryydrq9lrHEjuB1/NH1bu
ql6XV9OXxXfHmDrd3Q+7R+ikx6pA19fKV73ZmAcc8rDgAvyiqdheLEpyxY5gXy9/CLCKKh+oCQpo
ao8TB4LY/AFrtBmCUh00FzUUlcDGXySTZNRKZQaY1pRRITK9qYqq2EZiasivqHM0nnHndw/JSxGN
NX6C/OA24SfzgqDpc30qFCaHSAOUG5Xs1BiFO3BAt9hGPRCUJmWgVxLfe1QczkNSKPiRqY1H16Uy
0a+bVhaeOGX9XWSXSPApTEaOj1ayFbnKGYwung/ycmY4X6O5WBP6SDXdkEYoi4MPUEBN3XcILnjt
0T9nvgJACcV1DHMbbl9x5qnX2B1FoWi0URF71uSQUYywgsBSYSFdQLc9crr81YP4plZyvHpDz3rY
OnH4fNLTsikTIc5OZftngNQ/mGsE/opiodtBjRCZAQOIE8xf+ZMtAZfmX+uh/r3iHvz9F17vHICy
jigzcZWi4xFHpGPe98g0NVGtCiJNjhM+Xkn1nvU4qvMaxCM0Qn1GMvWl6ps5ogP+TqsINEnOAbzO
HpPUBWPWBHaaS8Kbuc27+Dm1moAbDVAqK6fWhbbfWmpcWyaEyr0PiRs0KDQV9Apy8e4XVw9b5r+h
DdNlDgNaioZGs5qu8AfoCKhOj2d8nN6Eb0uMSA04FmFrzvBXY1k0CYJEbky59EvrSXsbyz/Pw6wA
RTMdHXiNtW3UxvtejZAk1UTsEzl6XNap8pu8ZSfLe59rrM+oAX3UXiBLHO5EBJTEi27b6UQhxEO7
XHclikEY9QfO3ZjzZ6uumPdAiBvTcONVK54n7YnzNxgcjD1rHE00dmRsjTqvLMdWVmh9tTdylPxy
QAZUFs1cHAH1uwv9wBiiVjgv12HnMUJTMGokNXcX4RsSXAOnLpFyKeJfRx3ril7F02uDrJNQuMrm
OQA+Z83ixWz/wo+EXIMD80I7RAG1TeNAiEUNLABYENRqORlvub4C2j3pzP3jpriW68PiqntqEoY5
vjFs33Ia9TCbbooCsKwCpQefPXkd0uJsWvlhIjxdMh8W9+9E0WHrME8kr/yRa6iVgzcIfUxd11MT
59negeUzqdPrkSBXquJpj8Vf5B3glcA1RRkkilqtBTmPTpvNbtp0hqPHY1zmfHqh3KbT9Yec0RBK
fEnGH2TMbdJ/u/SrDm3N9aX/vmzbnZwgxleVoWmzI1/fr8Lba7sfWJlgCAYvqciQCQ6ePDV/s7on
cM4IkzhFtHEp3uhSV1vFCA1X/Z7ixxt03/xp2O1glr3uIYT/7m47Pc1qQ+sXuC49aI9ydtk0RTHy
2EPJFyCmrd0sQ+zS4rGdMuJtQBuMq5YUv2x1zehXPPS4dV2qew740bqYr9zeQeNVS23hwVg1DhoL
SOuCkoyPkTGuktAk9G2vn1JsYjZ9Tqurzgyar/zfQ8oO6+x/NhEWMy2OsQZPkJE6pLyYzjpknRxf
ptfbCMZCG7nU1p6JOiXpWmWwgrq0U/22O0YHrkFC+NbyU17iy45/32OcdcFPEdjnCRjghiOSDIIi
cWsVZYnecgHHN6nSrNdKJsCsq/gEfJZKRtokD2fltyLmNiegFERay1RkjkVitewzXGsPS0wcKlNZ
ggHEjA43E5UKkAniX1wgzt5OuUADMHh/1lH3X5NgH4bEr58cwRhtsoAdUO3+nh80+LnWR7M7/TLV
pMTwORHHNT0i5LmRAlYOJNe7j+w4Hv2yGUbRDjVatIoxJTNYV3l/NHVPXj+C2rSK5wehh/8pGipR
g3W4bHmeL/cpFYWVDusIxV5cEPoeFSUjGq7ePJUMKN1WoDSgOhLkUmVgLKI10iTAVJMFnn0cMSgn
vsmuodzaqPjNoSvK52ESgeRg1slvdtzDcgiSMuLc3fI2lzDN0zL3Dcg98t24dUxKNaHlpaH8pD80
+a1q6k6BeZdJD1JzEVz89yun4n6M691n17nTNR24PG7Q10m2JBvyMWJIAKANtHPnOIR/3mIp9/BK
gAB4y1Qrm9m4DUKj1XjoICGDUPCMC6e8bH0/x+zJp1cORil9JMrxrTJKZrZN4CpVXzxKFzWkbP3V
CfaDCGw8e/xw5ZioG97Rz08kULrWviV98zbvatDJ3hG72M4myRw/b7VAndARCJF2L0SiMm+u3CT3
2dM3y9tQPgPAeG//KsIK+3t8XFbmxyoQHFU8xJIv3SiWmM6rdLI2kad7VYADCkQw26JlqTdLlySv
GukozUAnMFi/VBgF4NDoa3qb86ve9D4XNSFgMCIP0WliyBAQxALctjPDIE4wyiNh1zkSnF7+ZtPg
+dIz0MrppDncSRBQyDAy2qqlySX0AsgAi1p8bvT/s/F29ricDamXocYwg3CSzC3e+pMWNJ4DNtDG
+/SVFS3YV2BIG2etPyn6+CR6yGAucb68D6rT6LEh/sQaxAL89unRjQcEL8svF0sM1K+LHWIG1VIJ
sMIXJMsc435fhFe0Qq1YINgtJc5vF2UuNMKJEVsNeD5ZGiCFpGUqUTdB1qJSDCf3H9cOcKUWhYJ9
XPNn6p2aYUVvzryPNOm1kSxBo2WQNqomCMPTLTNuHXAT25OH83NXnzkK1voz2WVqxgrWl2CdFZVT
kkYI7JntC4Vl/BeczcR+Jr1RgKrJhMshF4W1amNNtEMx++bSkGqsBdpKLcZ7f1L5bUxL66qjJYtC
aAvBNAKM2GirPJyd5JdFDdEpIEt9jo5mWQhzUDDOzRBI8nszJZiZ8UU9lrl1jNGdlTvM8MUi6+/s
hihBXgMFd/GJrLGgCQaNFsrO1/Ayx0DRrXkgGkzX0tV9vqPRZXGnbPRKhqQDobPP4b34JOZomckL
E3qlGWW3gMRGZKBaVLZeAeV4Q5lYOBzP2qGMVex3CyiI9ZaNCJQjVgwrSU32Pi33JotNvzafcW4i
yUB90G8PG23TNQ55fDdTj2qIbWlprltOB609sERY6Ef+tSZqGzr3WoLYvKZQc9J1OL9dtZd0Dxbf
xcWG2aQlxtZhKLf2kfc4KoQxbsAR9LdT/0gHVnYxHdeXxs1NxeLtASpw82n2d3eLEyLlOETBa6XW
kAKDkX5MpToHWU3ISZpiex+NHsXBry9+OD31ZGOa5xjc7QlrJrDEZqozkKFHmwHZfFxgkKG9J67m
7kofnUPZ8yYKX2TkVHAV+XRqraAXvFnhMqEmxtHdmw5AKVutSkGlQPl5IBXyVpjz3RiXVrTILy3B
P5NOw0ehGAss2MyaYOr6R23AUzvawfG5Fif2NNcl/zNOUcLD7NKrcU52oG9nrtHdf5oHsseCWvA7
2zY98S0eAk+m3gEMKtzjoFDoJGfWNaVbMlS3SOoh9fHcrdYlZed5K0bLmhjh7URoVRrOItmKGW2Z
y5suOvVCLjqyKB67Ax9bfze96DShKpix3bH06NBq0OBuWc6xTZ7X7aU2vNQN6wbfmE9HMbvJI3uL
OlJkur1Yxy/hSVQlKRROhAqPgwWwx67X3kyoVRZsstbENcHCNOv82X6HOvXP8UmUi1vg+t5cFIr5
aJhkfwe3g30cTxm4GF/I893SEan9PRbruJPQYH/ezzs/niVjw/XPD0TPEnQy4wnBYVuVSxIO6OS7
lEP98+8x/Y8f0P6w50PiF1WIpjwpRj9zKqD9ZILxETtdrzAEGm6O0REP2jahGswbo5VwNKnnKAPd
M/u/gwIEFuvV5q0GbT/RKG4sJSQiiO4DYNGu2B//ZuxT4sC8Siuhf/BfScVaTUzbcJ5XfMaB+CKq
/wmEe8JwCpz906ZBnnmZEDNoH2ESvVFJFakE5OId0Ova64CXsMK2vzBn83XAcqs2rSojsrfDhbUx
grpeH+HUjrGwAOwdHukZ2xG1QUZCu6yYLqoNfwzL1868CW2BjPI8FvGrKU44XIAz9RfUgsr+Izpn
E7V5NLqa2tFXRmMViV5glm16Zkk0wXwJ2Wj8w0xifPDeey1h7Jv6NkANMB2p9tho2l3vwgAWuVP7
ncbOMVEl9eCITdePjrpppr72y7TR1Yb8ydMkDHQ9QeDFJhQ5vLLfAGCJExsaSBb4CnFoSmRxv3hk
L1+74hNJvWPuklezrLtBjtsi2zKzvBO+oAgJYZ29Bacp51rsjA4LWfj7n4FR0sezCJ6dTIVtEP16
Y+L697DBcbiCiQMYY2FC4BZttmiAxAUVHmOlHcnPnXn2wZTzl1iQBDtbwySfUNhOT77l1o4hLPv1
9oA0moHjPGbR0UBzjiJolAlpqDkvKPgBAk3jXD6guq14n7G69MtYUPcT/B6/EGsBMbeIzYTj9dsC
TcnNXurEOILNbX7VFwAA2UO3BKOmNSk0w6/ZiV5/YdKUibjFuFKnikQ6Rp8HBT43x3zqCcIEJG9O
gIUgRcqdVEJskTSyoHI1PXCtxXjTt3QPSF773D94pj8onon+zpLEvpG62R36i7U90vetVhhr6zaU
ROX148U52IeSYJn3X+7i/5SrRxaxIPs/WR61pjf+LlZ7g25gWLExiebfOYnPcWehXAtPhNYBUYgs
RtmPhhtO8yGOFFJUnInolrsjOG0sxOe1d3kq4wihLjJzCKwELsoBU9x1ORReR1CfZnHGJEnH4qma
e2yni+K5vmqxGZGljf2p9vPQDACm4266SjJmyFxhF2DY2ANhG2uLxnK/AYGRvEsIYaKwv8F0Q3ZN
qLaX9fcpDxH55dfzTvSKprFBFhBEyW/LWEsunj9Uek7VITY5p5Vl/G0NQqoaCGLTt5eIyjd4tTL3
86Az3kdpxm/FatfJcT7oKoOxCJr0xk961F+4yd5N/vdNLsCFdlF8tfAZkvc33iAog8nSMUK7HtEu
3w3/Zm0ESwEI2O5d8VdXXIvY/ZWXD5LDfkMnSbIBIJNEzlrCO3M2EC9najKsAuS6/FrWwTMNR/8z
CQJnCV3TE/2UTVLglVWskRthDdxLZG8m3jTEq4+3cW2BBlIEZn+k+hwSzprrP/KiY74n1H32cBAv
A5wRdwGahyju+Dd8GljARnfkCSRM5jvAJnHebyWuPPXhvrmHQIaOyf000jFk/0nA1Ihac4PVrFy3
TG2a8H7RzxHE0dNW7XE57mRTtySzFpM9ZKyRqvw+OCUjnSrmeTPnbg/JkZZk24ydtuGc8vbkrkTP
shtuR5U7PkAuOJ4qpBVavX/MrhA2sEit2chWNxSYiQ3PxCi22zgbLQzCLXnrO3EJQ/S5Jey3trP3
I22wRKsySCDPt5fF6m46PE1LuaQH75yBLA0mZFBvstM4hXpX7837VK8dxhk/q3qvoWI7WyYjP3Nw
2xQY5nbXgwPQ3D0EuaZgVsWPE5OIvOvmp5plqCbXiXMN/uAYG3Eg19sijOkKfyiajEjttozdHvG9
HVPkHWEn2ZutAfTPLq3CA2h8DKijYEeYH0ord9wXsXGlEfTGqxZ1B0MT6nr0yiPS+3ajwW2ECsN2
sHxqMLMOrEvDcWW3UP7oq0AaXQbJopTgC3yo508ngS5Lcxv5lypS5XyovlPefniBZWWb72ZpwPF2
bKQCnCdY4ZFGqZNn77xKGC+XdNrsB5C6n94lNOYqod4jYndZe7kCoaL4EQhfvH8xmP7l8DpB92i/
w0qURf5mP3WyBDmx5Ep0fHtimyxym1DggKr0PzMvttrWrYcJJ6Gfz12vjjpp4Pv/vSN3jt1PRayH
VqfTO1SMrsh0TDFaZJZr25t48FxQD2QsBfm00QGxDSz0I+b9EwqPmGiXeWsTf0wHSdv2Dy1uhLV4
Kd7EnJaP5FdYtduVuI58oNJYYgT6TNuC6vpM/DSbd80NRa1ISG5fMiIsq5/+MD4T3AwxZxUY1l6/
rno5s8TskRNopwK493l19gkmXKpZo2nEOvlOVwMJhLMdtByMPYpRt62dKiZnCHjiktTrV2DnWBoU
OD8b9U2/Rfwv+QY0DeUZxG21JpuFIN+eNGtulkRkqiqeH0sl2xVcEGFp7vmhJ19H3RNcuWLs+qRi
qTeq6l6lIXLIZm/B0/BidiYF6HTEoOj3cSJwtMpunvCrfQxkV4uUUyla5T/i/np02N4C1Tc7L2rH
wuYwoVISP4UohUDKGx5sGl3CFKoAB3+ZPC3lQawmUEVFrtjp5A2Zhxt644xNm5zE94wiVAYiW0BR
3iA58tdF4rLw21xl/fOCg9nYba1Ro9nGriu0DjNmMPAmYHq7jsBMk/xMJtTNDG1Pde6UsqX0zXxO
zq4X1dh6Kyvh1jbP8KtnXA+Gr7TW6HgYCfIG00uisT/dB98uUSSgbYcZtHcKQ8dkzSLPGUcKhA+k
l0vWef2DI+KOTtEFQR3xNl42SgYK4t8JcvbhKxjZWpAFgIe4t0IdAisX4lbhTRHlh9OA4GpSl4Hn
8kC50fuRQb4aHTG59Istl/wm9N/+rO2YF8pFW35+l3GcG6O5hKpPtFOoQ7p+bw224Q84Gx6H6dyV
g4+g8SIgJTwNbd7rKfsyNQm7/t0GccSlJUiXW0SDhxT9kSbZqwLdbjo+9sWGoNMbQsP1B3w349eb
TBibpjC4eD+QiO8baeJzhumpHVZTBDB6LpNnZS1URzF6eT658UKkbxDjO9MPvYiIWED/SLhbIadM
VPcB7dzARqw2hVRsyVvZV0MpWw4G508fMaCeIGAmu2n/Jq8HZRd767dmYt88Uaga69emVqP2wv9R
FnjXJIotXZwfgIY5ufxaTnMGTNs9y7IjM6qZPWqZHnuG2sVJw347EflTZH5zJ2WrLZE/syDvFeFb
BinbeIK91brvmvXyQOfU1u6b7f/MlBorSe0lqEY8KYJNlrUC9PrO0IEiqwGph3LLe19mhB+6VV+w
VXJGG5/+XE++DV42Ap9Sj0/FI6g7dfDWz1tQE7t/Q8X3NP0poLiujkXbaRO/3ZJsF3iwcmEbt/TH
8BN6JQxtOi9bDeLEeTzCwEgz9kTaq9sRg6QnEr7nbekthCZsDbhFQ7VRmxrWrzAhorPg1FT2KzH8
s/+Zvr9hZQXJeRep8nGfhSq7ZU3hn7kjr/WL3aPOBbDoajsbSDWYvdD8aV+r4ZpQCpT6fO4lmUax
70XfjnJ4pM8vaykIoNDFOmm7Cl/6OI0S6q4Xr5QJTULG9qZsu8lAyq2C6pmfr/steU4EzNW+2cJe
EWu5joPojk7dScyrE6UxTLeONnUb1f+hKXrdmYuIWPzoiRyDo1zk2pvMKBp/sr4wh1s/qF9PNlB/
B5UCtfGfBYDHLIUYiXXIJiOPqt6FkKoA18A1PCJ368p1/qghSvjiuRxmft0lYVExJaLOKHcEfpE5
Sx5rs4QltSW4W1z92ZSKcaq+XFZlIqhP5K2Pi5RBwYIxpk2VqX7KZwVGeXufGJo9OlL7b0Bgy+3r
mViAxoFjge6Sjmkh8KN7oUl+1PI2tSDWmqg0ejXDLjzxmpaPa6xfipbMEBowIexhnafOJZZFWzTo
N6gy93e1HIW44r6IZmmYDGkDaOy5Vcw9jHaK2zNUlzOU2x0GcM5gPwwkD3c6CKtxdXCUhmawXsHc
uGn7yGCYz7YGIiuCe/dAgSUnRJAxUL4wKsHod/o1RPhd3e19D1dvL/wgl6iSgKKnyKroijxGo97J
+62TkSJ17/4bnZQS6U22uzDKibI1x41r8y8JyL/ZO0+rNndNBXupiovTniDvgTvYfdyUnhuIo2bG
4O3b26XosehaKmr7NVtPkf6VyXQJLoERW07PvFj5ysa4/93LN67Irk06OjnOEhXcLZgHPZCLoEsa
RWabdIA2doydX8k9UWjJmMphkUUyAhL/f5sp6O3+xmvpt2F+7xIoVK5uJyua6mWVCPmyrXCR5mQ/
DsE+JGP++GEI2gfd+QlJp4wKFhJAxmYMx171MOTus2rz1RqickB7lfoLV1ArBobaDec3HSWymvif
jPbzcygweh6nQ/8eMp98oYwQ9Kn8ss3nxcwRQBbijzDh7o4T5PtjLD17T1b3jyWFoV6cgRz4HEFK
ogGOqjHte5HVGfEmbYYvKp+tzazwBB2p8fWLwSuHqhAOm7XKFWdW2JWnVIU4hsWRFW7ypyE7bsht
XBgl+erccpj4HzNS5R4raoydc830yrDJDhbEDU5PrOFUDEarIivsGHNx3zce8ClttB4u/Tdf+pWd
XXxx53HtnJZH55CP31gptBl0aHAEIXkMurYT87UMzkGQopeDFd8jrVirxowbMFb1AJrJbdrwos5G
vluD5BV4iVkSjHblt/ot3FNfsJWYyZgU8/QObfgzzyNqbLiwRUlt8nxbVzHtGjCmpwPxUGKyH4A0
1y6yie+aoxCj15nJM0/AhuTevN2faUTpkP5czo+MkHrOX/1ak6kxyrHy2rWrqU9SylgWnUK2MAIR
LALO+74WVzlgTocsPdPxte/GMwEGfdKQQuu3T8Wn+M8+ArnWyXZ7/50YZ399uWmlJ+r6Pr+bXCFt
un0u+SMmFhJ7NmDdXeSfUOlZSxdnJW1k7VBGXEue+wreuRB3x4Oky3XIOc2kL2mtvELWRHivP14P
ooMXtdhzXuy+dfdWuzdFnHYp4BeUt4C4vj9mpXd+8erk90KM20AvMLuPYC4C3LGO8Mmy4eqnbVpo
LZFTkZryyo97qYuZdma5OmfARa0Qf5S4ILSk8807Gs8BZ0n5hJyxZx4rmzNpHp++1eTEe3UjcfRQ
DgCTaK1fgGPC3etMWAvd7nUFT5xOpCsAKHgn2F0wu4vkhTmiPHfgUzT9HhSp7RXEi42Ullqkz9yY
pDOzNafy0iR+YKQpwMmNqL7xdj9YUye2PXNViXX8kad2HrJ0wSwasfE3P3E0QM2ooRNBcosTNGzB
u0E/uNovTAnvcSpviB6xjA4p0477VPWXY+7IlCET5rFZYH1HqpFfLrmijn0ErlIGIbe4fLcXcwW8
g2p+15I/EU1nCQPF/jm8mRth3E1P9Fl21mfx5T6vcYixCk1x3A1Q/4HI7Y7WE9IS2Qv+7Zxqw+7v
GiLYZY7YR0QGzlXDwbnExmh3fqNfsmLZxfsel83umb7BWcOz4vP5X2s41o1ugFBAiqljjoHcF910
D2CU7LYCGCOKV5qmkDH/55wVA6qtAMPuN4kONc1IMVW/jNYZfJBxRkEiMNX/jZjgTCDzUu4+jrQH
2v/iXsgHR6UUCdqgVlqJNICHaPHGpd+wXSI+yHTqLgUsddyIzWHKchDlFH7xx/sG+IChiTUgW7Gb
D1MD+yGUVO+lgWx6I3IatsVYqsJUidc4gRLU1UizNc5SYzWssHTZ9CEMcjBK7wE844B36hE4c29N
IxSBo2BiaXYoHshVWLiREh0IN+VpO49FPKCoAt8r0gTJrf7z/QnaKWsLIwb/uIeDF08bbq2QWgN4
cOK8t3J3lxQT0eQeLJu62iErPZfIFpxRohghyXhzQ1isoGmSBQFvGvXT+ZFFQP5yqriyiMQCmgmP
5kSZKd66QJLcwU66Ci3+bTJIy69Uql8g8YN+nJ0bh2QF2MFAT/hPQFLwuDrS51cJZsSqWgRsZ8vp
JBhxlG0M2iuDSXiAJDXlPBBuA77VKwfXfRWfZD+N1NTWXzwctNQvOeXd1vpALrAHVU+gB4NI3Lbn
JrGRjNAZKF/fAtilXsOeNwSkLPtNTyZjt+NA/SROEfYUZPEBoajNhMz2Y+UV5gp3tRIfnKGbcrbm
m28Q9OCwLyX+UBwJB3NDfn0aaK9lzb4oPyc5bhZEqDG11jSP/ZnTL+fW0RMkJYy7Xn0bBL4Feijo
fBXGyfiwbXHg5PCwWePCrNndosOSRttXTq45Dmdnx48BOZeACi8sg84Ie5wdLizwV9FYOekwxeX0
lFq3cT3bXZwSVzjZyVcc3QuC1bY3eGZWosQ1SPLJ/DEd71Q5dp85MbUzaWQwvT8l1K9tQMeysGj7
AgkZ0xLbhU5d+NNTaIgOOdWY+cmzz29+YsjHBeQspglAtFCmT723oa/CvO48sEQZMiujWrWDNK3q
MlHpjiQdy9+WKTNZmNyMB60/KJUTtSuuCiwqduVDf4Imy9WfIBpwVmGcfivVers6N7SwJui3UEh4
ShXxQVYCxjq966P+SOSCvuZK75r1QQJIWKyKpjTFD4U0pFPyq4qcStK/iJg18aduY+I9LyZagm7b
fpu4ioT9JN0rvYbczceBTbyThgweA81If50qz6Pdgst0j6MNtL9FhhbwRKb4GfKy9gc9tzlkt+Wn
tNXg1jhQJ9I/6iAN+pT+54BDbIwOIYG0A4Cvg1EdLb30uT3KLe9JESmDfvHBZg3iGvpNpojhhby+
MWnXYqnzrQRDvMkxaW6VAkkXWCLY24NU+51B8v8C4gCTaQeB4aeAbcLHUO+OytlXwDWbqZ3dQ/77
GTjljVp2vWmYKGZaxCPGN+0FUroi0L0UylHw7BfC/8Q1432Ni2AXPiJZVLu4PZKuuukdWgtPWgob
p6kQ7xib+lfz/s2Q5V5lzJNpa79D5AJGgYQAYK6JAqB4as3T5tmxerrzhLEQei62J4raVL9/ucwv
s1+uoVmZGZdHGq51qNXKEVd7HoYCJtTdYgnDkHrXBya70vjmRS7EPh0UixFbtrmg1J45UiCgNz0V
k+CGK1imPBW5xaN1g64B39Sb2moy2s+s0IDAX71wI2eIYnldbEg9SwN8M0vA94V6EwxGbZhAYtAt
yRXQ8/k1RQoJtstfxwkflqa6/EZz0oVRWyYW9ndZX+X1LV7og7TOemQMNyGP06L9Qkch0pZPbp3D
Yv00drfeyX/pnYAWY4py8SPDOO/W1fpVLcGw/2zE280Moe0NfwPc5ITDo+fM1zRwqMCtgPeuYOW0
a08kr604cvn6fcvGrC9vbtkqDC9+lRbp50VpSasKpTYGzWaD/21o8jR7IPblPBJlL4rKFVRSTxon
ZUKAtXiiUbnRzXHkqLvwY8NYgdPTYgIznvo+96PHt/bVT99Q0PHOZT9WWViXOh4l/35QSlfwpaSo
3y8J1uZ4+HgMy584mVgJqk4wD/Oz3M2gtxAoWPh1zG46HXLHQumPNpeWHJWcI/tNUkZEaLiavnAt
K6Ib/DQ5a7o9YhdxAyaBEAdsif8ZeNsQwLWbPkBKtRLSOeN0JbH9vhkD0XocQiQ6Wd6bb+wd+d7R
rNBHKdl2EXKAzCVjXhm4IAVaJFOxWW9LQMrxonKsA+ubcYY37KXUWPArJSC1u/tlGTdZHdvJVcvF
MoB7vQaElIfoXZYZcI0AID+fvzy4oqb3u+R7GwhQNgZubE0FwAc9kNHURhnGVh9c2ahMRr78ONz5
HJkdPTThrxUNCK6Ht1RjGnu6PWR0+JPGldxF/pWN6dgiLWp91E/Oc3VrbDD0HNECe7/4wKBtDxjb
2o1bSrd12UoHVa9xpnEcwKHpX26VRM/WemhyCZzJcNxCPyqi013OI0i9tLOwv28ZnboV6EaeFU2Q
TF9eAU//JHXFfUybXwsXJVypCxjTWkoygJAYp+UFmxtWAjOm2YIrf6h6Ckjeb96bFn7RV9fQ2AW5
7lXfYA2X7aY0nCfYXjpXzJACiI9AuVm3eJTd+Dl9LC+CrLxT31S/o2GR9GmDAh88+aQ7NJ/CQEXv
mPS0FVq6zQjJzbld+e7eddfwYG25FYGfcwT+NXaVpZxkYLz06q6ivyrCl/2D/j3/AWyBXNGRCIne
gXyFArWO1fW8WoOjXf9SMEaHFd1ykol32bXzTnqV6VQyJ18Ckn1EiJYmZLeD0QK8nr0W53AbPC03
7s57M5okwox0xbcBPLERkBGgvL/5f6Dc2cm8B85yTHetEejz3fb2ZqXSvvmEaqvX+6196aV3p9ap
tpcbEipj4GmAkjM5MX5VpEscQIVqcnVsOzxsoDZuI9z7x/ZH7KY5X0Pi2aqa/ENzBk/bc/vIuh0h
C0kcSNWXKOnlYGASJiPuFfAFJ5wWfcYCPW7i/CWc6oV8EMRGfqnBQr4FsXvamNnYXSbiUpWt1Ile
dkerLQ4t/qzWDL75yMMVb5FF/lgVxhjUbAer5ILY+TiQisS5MU4hcyjJWplZ9ZDqx1aKUDunQL9j
ryt/YsOSdSvjTaf7caEC/kYhpd0dr12Gn4iIOcUmJWM1L/wWJ6Gvot9r9QplV5YTfJjZy7oDyNU/
yh1NpTe6mQ2Obxhrv9zKsT+Ub2Gyhi2cqYEKEYMJmTfRNtVdTPM7pK765X80Khvnbj4QOidjc/Ep
ZF1BVzDJftrPIF2wQs0JJahzaQCrI8I94lasK7Lwo9ak/o93nEP6SQ53uDo90CvuutKyDG4hlDmx
SmMk2qOHEnyWGxw+44aoimvr1snmVUQwEHSXf9Ba+XbzNctUB1h9z0yxIEX1QgIeE/wpbpcAHKXo
R7XsokFtjvBRuqIDYFMUXTeL3xZCmXUQe7Kl7LFBzPXSi+pfTqysPnR+Bj+VfEhvdQ8o1Hdw/+Dq
y165FYspcgWcf2JEA3q5v8QKkJud2egoU9AvvmMabdGpdrg2+/1RwBidJg9/YcCJ/Y4QEBt5nQe7
0jaHcMv7YXhSshuAC6bgiF2eH7bt2ycZjOl73gNWiisOpVAjOiP4pjyorWyfxqwR3veiEzIBZCFB
O+t4aJ0ikx5JNAt02bvGQMKjweAwIUM1/RWAyslWyU1I+c9xoUvdUk41a4NBMJDsY524B58MYv/o
uAvQPDV3PfaGTlMPUpYhiBy2fAY4ro7Vlksx9U2zgtBGDswuoMn85fxifqgyebM18SS/fF/ZYyOJ
RKwuUaAK1oxSoAy7Feuuyj84/mLy3rTgV+Tr95BzoO/oy7N6eaRz4z8BhcbkL1rSqcaysMmAFQJj
x8W3+fRnQPx99J6hbwGv6TKyh1dylrYgRTQn37Wdo4Ht0X4aON7PXSlzc2vxbxHIDTceVQZf+PZx
oo8qEdP/E+ux3CSmVvWvZa2U9og/KOxBTwbnawJc4YqkAyDYB4NaEm2f6xwh+UUy718UHlUU2coI
XelJbOkjN/vheUKlQrmN3zORgj1KABgvJ8d+zr2sQBx+JKPy+Gncvwhfex/SveJSYJLIW7a92ICb
sZ+UjQHgqxfv7WiDrW4Fl/HTeVfehmyTfjQqa8Yfdn2ED49TJYpOdPlESWsO5/3UaZjnbVGx+XWV
WcrTbPbBL9H2XZf1moU3OQ5nW8rEwrwZg5mMPl4KAmSUVwuzfeRsekJnsn90haSIS0gdi2b7eFNO
PjbiFzzsIlsF0zfcVT++f27FObh3P6zKWZWL4qi7toJdhkBLJgE8jF/PpmjK4OPN8dTUcd5KMAUq
s3olEU99WZ11e6UCfEwdOPbHOi6HgRdWOd4w1zj8AqbnT4/2eW6hUqPWzPMFy4k7jB/h8nUVJ5se
/Pm7YlV3fX6zg54DjUxlrlMnU1T4dsN9QPhKtDN1tMLAWwSY0aId9gM3zUqZh4VOZdduOUHPqOpO
btXl9xZabiKtPQdr5ruy+8pJmEgAnoXelyskBBnE6I40ezxCBfp2yIXFYfCNae07iopzYl/iBIt5
+USrRHmtX5P7OdADyIz8iLasoVYK4LBTyI3/BaEl7UyOakmevUDabuUzrmGBtrHMshCr19dq6S4o
l3rqsn/N3tFhVhBehYGa4qBLSvXcDk6heXo7AHU5Qou1K0Q8gucbfZ1t/9+s92GSvf48RMncjgJ+
cLB1t6T4wm4Wi0BoEziNejt09667Ba62uT13XfaopLiEC39YuvZBqbsOMOyGpP4jJHwFMCz3VQrM
18i8Qi2LNwjHkFNsLz0oihew080uqEItbLjNUPKVKa+jJiGUOxMIUf56aGLYJ0i6yMfa5czBbU0f
uuKLCj0Vgau9QxuXGVu8Khqoi1OMGPdsH1qVWY3mX27zpdsHWcNk61/gSjO3yHwapquHhrpABXlw
rWjKTXZ7QBvq+f6I4k/kiZdtsdeJrk2XcMm3EPtS3xoxHWvkWJbGdel1+hMuTD3sErETFlsrDs53
1PFi9udIKKEUe3KSp5n0XKDEuQ+yBa6SiAw1tLZ7RTSyWq2wlAOZfq+FSN43UYv/J4hw+DRN/945
tqP9pLEA33McigaNJW4heze6Szevl6rbVGD+tntV18cbDyV7vh0Ej+zvIcvwX6z/tPBZoc+Xggix
P+BIYXr3GqyIVVpiiPAe0gaM6AQzKvPkYx7Q9gTrvztT407SXLwZoWg59uihMbkCDMHEOoxc2/iU
Ejynu2v97g1THGPFXRmSreiKIH2vyIcvJ+zjBonZp2NeloyY3i9UmVo9asRVer8vmanTM6XbzW3O
tTTks3ZSWlZ0pE/dSbVK0jzAiaYJ9zSiUEnP8GlSra/iokf+lETrD52DJp9Ht3l+rkdInP8G8j1D
kwfY457ID/8poW1Gqd5MbPx4TpZkzw9hdDUAlSU5+WzFjDRETiF+mkssTE9H5Xb4O1p5yj9w60m1
acR+jc3FyTVolajTJtmlv+cso1wLgFi+cT1sbpppGDnR/AxMzNUudwwqSL5eVk3acVgenzTTbHhA
AeAjX9QzPo4hb6d1ljG0SSsn3KxNvjsnToAbp9LcFsLGOD6fTMq33JOX0VEc38n908FvpAWZWSOW
rV1ONpuc62hheEJyVup+8w6fnRr4nHXOsa8HcZnSO64pkkrLV884NHpun8JmffQSgB0788Sx50jI
59vBt0Gy6Ic7cb7ik2BUIWWZ0TFa03MtmqPfoS8cAEkX71wLul0DS2Ax8c16E6Q6MzB5tyZT4uLA
HQgFGOhdIFaaw5ILlWQhhVCGtw1j8tBKDhFNSvpIMtF/sQkF62rm9u1cG/+YG6Ul7znHRKrZPEjX
rfZmivGkVAZHKgojtIqI+qMqq/HTW5N9Yn+sB2s72IDgDL+3QCgkDDMpPqbrQf7tLtZWbCAxfSVP
c5WPJFq4hxmW5agzsGs/3XlF8N7f3zBGuDNEHq9LQXomz6v3mabLSdEid3r6bgut1W58dwdrEnPH
ZlyAAmdAdZKLZemGWSG8zEQQI3NT77dmHzpU3Zbbsi9bv0mf3vBPImIz3wKvb9mZGtiB6Wj5tB6Q
Cinvlf04UQIGJQ61BYuFjuiwV9pN+az/G2keUqt74DDdYjDQ2Ryb1Z8OfYxI0Bj2ofQrGSHDi7ln
nUzttdAmrhDREOZwy1LbzKU0DyJ1njezwkwTfzMIGJME56yahxQ1/uQKSCUKRNoTNh5f7txBdabO
lp63ImM0pVqMZoULxrK6u08P1YCaEX/oNJpGQGeofkPQHoIvl4Iqlk//iWms/gvgaA4bTShTq7Rr
G8vDDQMdIudM3uWlQuige5UV4zcSolgLQpBGsNF61d51Mw0zxXMeASB2BD6TBuwYBHPNWr0x5K/E
oMRigoRgZHyFt6223lz0reS1KnGibyfJzKb3PxiFguQjiR3sV3/W/kHrxryn0bF0O2mymq3TtSRo
H16mN9cnlyJXbReBNt9lNkMO29c0vpmCEOpR+dYqqggaHTCoMNdm862+AEEgNBBdpy3peEFu4/C2
1uO7Th2pF3N5yH7TJeMUuCpE0MGcYymtB/kwbXBAcGC2UmwTSA1EAIp1eM3N2ASZNivqth1VR4rc
7wnGYFIITj+zdibefp9OuOFAuLr3BvmHRNUlQ7+p3OWq0fxqrVD5GtXQx9wR6fYCInaVcjJWvAxg
Bc/w6eemUcq5HQi77Zsec/P0su6USYQpp27+OYTM2/DnRW5yZreoZpKLsVk/RtIFwrupRMMEgjNX
wm0FrwkuBOrY9+vc7Xv8tptxf6nnYMmJeOnZsXVXFyVDAA1y+wbWf37cKjHFibEpzK7DCPazy8p4
/lTzj3ZVizxI5uOiHTdr4DOtR+gNeIMPxtkGnO94SngbkFwgGvF2hpSrmFNp1oqcLfvcQydp89fL
VtgGTQ8eBW3QuJaeXwP2xiTDzwNrXG7zZKHpW8dBYX/nJvFsIVLAWyyWIbbnXenrcx0/EDIGajaG
kKbe7zm7M+7ZcYTIvWwgoRPaHDYN2mMLWWV3Fp0HjSyoeBcHzXSC+Ma0Cw36kbTPMLbxX+I93n7g
a9Hd5RVq5aQlGUJn3unC1mvjijsf8xPXBMKcVBDJPN75P+CBXSmXN+u7LkYF6/eWuU0oBzG1sfWu
pP9xJGsaoJAD8YQZXfVsAV3vRmHbqi5xW/EgZtdmxjxPhkKfsgF/IOklxBIsnZybvQ2R8Ly+eFP9
S/1iouCuRWdMTWhBTwttZ3xR7pE/OPdGe5nBX+lgKFYpqls9MmkXctJPR2LlK8wj8u4tVF9UrN1b
ThNlbBRMV3L1SEnaTMOGREg+n2H8GS6Psq9jIw87dN7aicHgFfRSq+7SuakHz5WwDWRaWv+jZIG5
razIEDpW8XNq8P4zjwUW0fWzoLsHfg60FvWs/6Y0FwrfeRu7XmWM7nRJu+fA4g/3ITkktW9KBc+7
SZncoDLKC2uJZ+H6iWYuQT3wXgzHhJLHZEaNz/2bWGOVV1KZEiaOuBolt15UB8dQ757hg43Gbai2
YupLf1jBoLU9oJ8vkTYhsZ8bM1IjDhj6BQpOMmub9JNYQT02QuSe1gTSENYG7eYcwpQULkyvpFsj
1BVS6jTlajASGJ7JBQvNkniO2XGIejHuHtze0mLXrPsJ5a1V8UWc34NDMRXSI99Liw/m8rmb9L5Q
FwwbRpCcvXy8K5Ko2/ZiUhUN81iQGOtNSx2EA+HTMCctZgq8tFlwLsOyp2tbIvPvSSwHphTF11mb
hxiscZIGeKue1/OgKW4tTDne+dEioxxBMoCV/hORMjBvH2talSIa7iAXWtdDH+Q0rkaac37Sj8nk
JElczIKS24SesU0UhLtnMtqgRy9uHAKYb/oiY5IKRvuqVp8hYbzNvy3oDYOsdl7WFsrzSFMqJk/0
j1ySZPWChlxLBnDsd69jPKbiHnGN9FAbHN9X15rOeB1ypOBmmb1aRIHe//cJdqtzTXQu0GpJwUSR
jAUPqctwvZdzNnyBHWTAYHu4JU79gJHzOighwZjdf8bkXZacZZG2bkI0jL6PbJKXda6vGorpSHtW
pixgqVIkkTIt6I4vSYGla7JSYdKVdZ4r3GUX+HYkrkr/kChfsl6dVjjWluYhJ57kqnqi0JYlBeId
U/2S0z/etGy4/RezVqbKn2gutrd6jpxHGyYKXo7Q+l6VoMBUr31NfaTFFr2B9ZhnctSKtt6lKL9r
R5FUwx76+kbP+KlAA+/PvDuF6Oi4vN/q9EOSG9ZYFBefjoNgaUG1uGGHB66FHkaml9lx9b9RMmE4
4UM5n8itd0YsHWdQ7IyMrK+CPOct4bxVYXRRDmnX+96sGHPIBtNDvEtriqRz2jEWGCKuZ4bMXKvE
4SiNZaaA5tsRVYPw60m/YrVDjcR8tJ9zFcYkknQTdukKU9B9gk7I3v6JUKjrVDG4q809bQec60a9
xDm04L+SESnWSjDA1Q85Sk86ElpMEi0kXlqo4EYiinE0pvpwKL2JX12mqvDLbSkxNV+PO9wzrH1u
HCsHCaKXnxQzmjcGKqFnen+oCGxaAsD2a+rJeuQSpKkWmkvR8LVmKwtMoTWCvaqyNKt/nsP5fROJ
AlTZOY0N1mAQ46LgOGgzihJfP+i0HH4mqTNKBT5Dg5dS4Yh16nPuE8vSe86h5I6dcZxY3cMikGVr
vY3rgJQ7zgb1XpRMFSk39Yf/cENPEiO/iyvNsC2GBpvIkDzMPbbV2oz9iLDtRuitJpL8aC3sJerZ
QxYkvROVp4cYrTRKZXTJAz4/DRRoaAaeJ1/pEe4Ffb/lAACcfMe6WO+qPLbUThaWSdMiARSylpgx
fDAKnZsKqJuwhdmdZfX1oJ4EugzOgQCu2al16UaJiFb0MdvSi4JePu2TVa/M0WG751K9a3Q7Numg
ZFw2Mz42NPhamDfJoEiXQw2/1UEF/zxbadYMSiIs6fhCUOwbEKzey3PZQYBxr+D4CHn8dokSlKvi
e9aXzVIX00Y19/xcJtC/aqxy+PKTWPjE7pDDjCVZ/uCpqWQ4NAHsc8Ye9gmforSofcb19VJXJFE0
GAD05blaRSUii3ygbf3fa2A4mpvYufL9bEv8iuSeIzSClzw3akDUVh4B/WZ4IUu9M4Mu9c13K2HE
4ssQJWArdZAEzE2CjD2YQjKkWAN+zTf7Jor14rS2Faqev3eheho69tLwZjJhOMAcBoBmYwW90YyT
TjWeugQJTMB3aq44LCNrkqFuPeX0EzAFoyOfDsYhPubxQXY/Ta+aztOuDG+dh+cYRvkWEsgWicx0
0iQVjZg+QjJZ/zJviQHsiuRXvv07v6vnJ2f+1aYGAgVr69VWE11lMjELng460DNueDLtYrbx0UdJ
JHZttXaBoUsUQQysF1tUgkBlv6dwBo4PHK38YKvctUbnv3+Jp2PALovahJgfHYG6yUBDOWAkFIjP
gWRRN3Lk6gvWy//FjNvzGeQ5HZGW8LPhCWHygPyUviTJ3NcKSNrcdD+/xyhFaPe8da28kSwmOXPy
zNDg8pLd8HLd3Jkr3i+ptdiGUjbwTr0Gn4+lZorqJCk50h3bBUh/oW4HqrPny9MHIipHFh82EXP6
lRW//rv4l0nZI0Nolu50EA9mUUBtIrSBuRuk5BPuYH3D4uytpp/jgdIwppi8YNBZJ6CmG/kUWYEi
xGs/fvrVK1m5r1ce+vvZVjdrldJWmfDViCxA6UuGhks4U0sQTyEVTl8jsDOviMVfnLBwUn+1Kc67
vYnWMxeUDMc6BL4H4chclj5mvrKQiap7k2Z6QsOy2vonHPxMgJSGsqD/+9jzUCMEYP/59SpqXQ/+
i4Ieso06+RCASSezg14OTjpniZsuZe/vz0EuuhglUGYplppX/jQCPqRr6v40IKEE6zEaficveAwv
eWx3fCPqyBjkNIbPotYfvQIUET6kzQWW2fnHbDdwRKcuXBTQ3qjiIjJGd0icQ0VOPKukLHa4YLy8
I/670aQfywDHMdM3DdOud0KyyaL/zaRutrLpWR7ECILGdbj3+vjLmUsnAMFUQg39mJwOZzD5SeP6
crOt0eUVKGBYZhWolcT+Afywc6r2qAmC8PbPPsBRjApaAU7JPUdStWD1OoevhBDMPliIhGoXrdUW
4RxWWyf0GcP1ddd/Mn4DW9BaaqXCoSFELBVw5zeU9M8zKdTjjC9F4znOvtW6LEgjGkplfyWH2Wyj
fW/nZnHCNYDprnfJ0UAZOPFrzH/DWTLE0cmZ312R6s6QPHAGqcKg+F8QnlP7D0uuEKV6m+H4klPt
Hv6zwO1O0xMCD63y2AD2SgWmjgoxZ/2jCmcrQrG7Hl4qRF6vBg4q5OjnBb+QCTdppNlnWhPtYDrr
I7OspkCvZteJU2qh2v4lg/Rf9wyZqbUIVaBhbuq3AD3hhESY17rdAfSHd4c7QzwHB3abTYLlaG3A
qjQ0AwjKfTCUGmIHNl6doke25dcQEYCKwo5FTfWWSwQlJDTu66Qahh+uPJphfhL+0Fh+ugMQRQrm
3ycUoVfOqm0pRsT+OtlvNiumX9hO3782zc4MaoFKqNQcoaTaW21bXTQWX2H2thJ5d4hPlObg6vuE
i5f5aKE3yJwHiULN6yH6Tn6wflFfXJPl3xHQTORuFXjC0modzScGvs7ze1kg/mKuPuXflzDXuATf
OcLOAGA0dG4q9pVOovAPRq2pt4EqcSdHUGWoavZV9sb1+xGiqSeKfBJ3HHlMFpw8Sd0hoWUVPnAS
wgYC7AuPNsq0EAQbflwfW4PqtTEWgJx8pikV2EkVbunEVRuiac+eE40GIyH0x9H65vwUEa2OHElj
jm4KjcOOhr6Vhfay4cqSbkXFJ0e3W7jGRFg0EIecF1DXWGtpI9oK+TLI5QWMKUO+SXgu2KstCtnL
b8x9d1hKrs7i7ya/XywlOksoa9R9voadyvh3W44d6L8xcAxJ/bFONbIY+DtBx0QatCEgzrb0OFtM
Lb9pRDzTy1EYEZmqCd8D9jJd7IBw4mApNPZmI1Tt13hAOYggmYddsAIayj7R4y8CX9+6YrEwi0ps
zKqQLgJz2PTLsMynS7/0L7hb55fwidrG3VFuSI4UisLCCkpCgNQYUbJrzsjYRtJs8EbNtrYjV71e
ywkRAnrJn3oGrYjJ9p7WvjnGh0P5O7ZjhWmM1wnUDWA2l5I7+J27LQu5/B35gvCWkzfTc1DeqF5K
rQVvU5zfWG64m7DrWUbpZI5enKYApRjD0YCHRONXleoTBNInhPznMVKNbUmWXCM/8YBojvTSRAqt
wtZANd6MvQ6pB9TpEuIcijaMd7tXWDwgs3wVeXjuexh2f56ClzGwD1Mu+c5GVvLH/g00kUPKP/fB
WFzZAkeeKfy/o3Uc5mBET+hvSoSvNLMIAj5ZWZ6r6HQlqT2aLhoeTBMhSOCH2eqnhFkw+pEPfzuE
t34kk72K7RH1GSCvyDsB1BbxY1x7BYxXeZaXTLZTa0y5ZvNRWOzFWVliyuykbgGx4pK9nG8lL37m
S+zJt6+4v2sIoOZU0i6NA9EMQpyDpMpXFipj2k0w6LYLdhiCESkLiqqMH7MkK9sB3ue0iLXqo0yu
KYRo0MgcgFDjg1n2WeatacXlPN3Gy1/0FVxX+q8elP84ecgDlYMNeuFkcvc2cR4oR/KGSsODk0Up
Gjgo9jddNtnL8DoPRxTi6+dxedI0+J52X2r68IvLHqs6pdVOZLR5Qr4Dw3CUXsiywV11r8LOne4r
XGPB8hGLbKjuDj8gMtmQDbubWNFXuH+l7w4KRbYLVmKAQGYN20xucE6gJwiMbdPdoQTnjY8PXdtx
7aVajdshurITvjLTJtt0s0qzrFJeshHnIVHw0HMBy0a3Y2yJFvKbatxC0b4bPgis3diTUIgEDgeX
dIfNgqDbUs1mM9QCmI7Arc7dsILDqavrDwbFy8zFP8c/CgZFByC3bz4PDkSnQyelexQFhhnCnu74
0+U5/X3Fzodkupjk8G/3ZaTlG8nqTLtBjtuq5Vzj0vs6eMBz4NJfcbtj4+JHyfNRhlDsyD6iQcIs
yZ+9VktO//vKKbn2MfJymBDylzZLvtILzlulAPthAK57EFGdZN9v+SMGSyp82DYXXXqRH59HPxYl
Q1tQRmwlSb3Fskq0TJ50BepKGQPwAItDwfxpg6d1pSKOClg7MvrwRJoKcHgn5YQPGDwXbcMamDNQ
Py4Vl97O0eUzO4P0s/I4TY7equ0zmEPJ86YPKycxuZCWXVF1yMiHHpTUGOOZ5uObtMGGQ1TC0LsX
OqS9gXl19bDXVSW05ZCJnv1XSI8bSffGVkt0HQpzt2nBHRE9RtYi4B0mQfHRcFXv6+K61GL2CYG4
11zHNV8JtRdIAhpMQNn49nWqU4mw/+9Q0r9ekT/k7LkKG5wTVy6v1Kckh1V5C0FwciwHcK+FDj78
wNK+Zi7IFRPIDFDZYg1N2+8d+IztMwjS+kDfyCAItT/vOu8NLZfo4kWCKUCI9UXgnJZCxxr3pAIj
h0xBLVeEf3i/k6HiVQBUO9FeTlgYzipb8Mz90aL8F4YuWhdR6hLrOAxOQIo03SdNfXoxnaTu4ZZr
1QrYtA25mhQCI4afBRqq+E3vfVfQKrsV7fwzi7U8WL927cMfrDsfBMcauLUxd/LXUnhnBGSwIYZq
9bUGAg2b/Ys0/ReU2cXlV2QWQV5S/bqFwqEDmjHqn1EbL0HsXoXFx8VDjMLksEAEZAmaolH2lxCb
4UPjofea+Hv+y4td1jrWDdFIOS/P0D/IN1UX013xRYaiYMwo6fqMDmB1tEpXtmQ52SisWJXP6JAd
0ISyWU+9KltN38zMsCYt1DpR5N/9WVELZCTADywQpI1XUQsZHf/OyP1/TXZxjsRiEuPZKrxGIWkQ
ezGwSqAvaXSfUyldeSSnTK/XaAbajN5IYFQQH2frTGVXHpW0s4TYlGjr8YPyhD8sIGe/hGuAwN+b
JCkdDWK4IzWfAy1KTIVAHed8jDaPdVFzySO7FtUQuwT+4UBHp/YLEAvKScbgIYUV5wDp3kt2cqaQ
iURm0c2y/S28HFygSMnsHQUVee0XqCwlk7r3uFQpCfyH6HZzu4YLz9xtAbmZg1G5VrL0Lvxtfgte
ZdNZ4NdS7KCB1wqv9kzocfxWTBnbUScv+dVn98LF82rkT1XMrTxs6dOB61u3kgeSUOCF9xEHo4yi
bA5VO12MhXuYh7+ZY7FmiNabd9dv1UUfqEHKAJRn7MN71f9KDmmf0LjtxTHVf0kmaJaqp6LakLvt
1imVxIuIY0h4uy5VO3lpkJlliXppvTwCOEWJCy1nNosERerkG/fU4+Hjkhmz6D4I+plcIyC+RnPR
K1NQa65lAiHqH4va32+mfDazg3F0LXGOoNbxUcl0P4ULlsO/8Ieex1HMCtWO36Kv81ZDoyhOxCBh
NtFWGzr6xREIhMQbWk8+SiTejSJ/TQeuEXQRWIbjnapPXV7EYFLpuGIVSbB3kvGY1CarpHRMoDgf
2bHZcdWI1DuXhrLVSEZsAJbu8315A8iWWMeFVv1bloNIyTdlnAmRslCeetwiQDEalDtTFcXLw+Qh
PkNR6Txkj0zO8xnLtHqD06QSUOJqVswylKoE0d0ev2huFnmHohaHth/XSPFwbQ6w6QcSlnk/ZLH6
WtBYKWVRN9MATq7KlQ0gE5Yq2F6yC0joqsseBVO05VpAoz/DV7FGq3YXYrtvaRoqa47SKOrXGj4v
VdEk6nHk1ZYJE9CWZBJt41kFMvTXiW+8QvMxHSnD/edrC9rBt3f/u+yqORPhWx89d1lQ6VESUhr8
8FFlEaAay/fl65FZRpbXuT75QjhXj8J+NcmO51HSELbGhoyDzkm+qs1ET2KmO90jnWT+7QNmTzoJ
BhBuug46vkMiey9siCGCJqu+yE34ohCp8wwmLXgIS6hXlKdT29EJ9g181qI8bD6qHtwLkGj6fZEd
QDyYDVUANuDUxkLQ/6X0FIVHxaFV1uARQ8i2GoM1vMcj76jj5zCpRvUx1DPMaTdgHB0Z1m/AThkY
RO/v0DdhYCE/eY8GNYOn+TgumEq+BttOFhxpsLd+ckavDhbV+35MI28ygTznxTABxN4bQES9KAfR
lYSXizl2vUnC8pSM+5+lgEgOuUBiZ6u6Dt2Zr+ox9+/AheIVEOG6dQCLplXZrPyFxu+tq42uzn6g
1rb9ycfBb/qhlesDgiTJ9a/Dmbp9EPB3RHQHFG+1DWLSA/ubzEQwFb2PuddGJ0C8jDrgqYCx62kM
pquiHPofMI54MpFANboGU9j6hho3NxvVSFyHc5+u8+2e0DngySeaSrC4IeUKVYgM4+RFpXbjVBs5
Gg9ZRJmrd5dyf4nj6T5ll8DP+CM7KrAmA4zTV+/ca5Lcnbb2zEkhcNWZTcPZrjA4LdylB6qTrEhY
30r7xPtlDqQixTI8biDzuD3ItDxOqCc4u3hj+3/+TnmL2wMif3vw6cDeX0VUzQrstb9bchRLTPlQ
R625VWB9fqyboX5jJtFak7Lv57K1R97FrLPKEfuArLuxW50JzkmoqjhYmKt0i6DgTopKr6y8qnPU
u8PzJG8AZIBTbJUQxA/XBms78HruGpwXHI5en/rdza1Ayz5+kt22UU/Yczh0QC1ef8ePuoJqYF8l
+899TbuFf2GoMcD41n1UuqqZvkbRAi8UNFcusfbBv8yUGf5unNlOy9t+yNjk5PG77lw6Bv6SFo+8
i/x5PxBHCPJBO4pG3i8EZL+ncd8RhxDSeDDWOPGPez5cLhEAnwQ37g/WcZBG4dCanX3r+kcpQOf3
l6/lwUy5ESbNEafafhJuS3ftrtncxmbgiJq7xa3j94/1aGtBWo99HqsIea6xYmRlFoAoI1ClRUYQ
ecXagntE0PJM2UpAPIBrDiiq9lc+CR0cigdzU60WXM9ge75SLHlXS8Qyve4OHS8CcWDIzJmY/9wU
EFZD4bBr9X2rdbofH9TcyD3ObQ835iJT3/n0X/koOpvf6B+UXe2zEK8xb9rhGxXU05DD698j8VLz
URrTz8Cuc6bzqJIYM6zJAYhhZ67BfEqe6ocRFnz/ik+ANIUkjtE/XaoEnym8ybjG7/YinBnWpCtt
t+g9cUOZzzRDWfn1l9BSAYfP6UzihsMyz5obhmprOLIiDQ8A8fojqni475YuZKTM+3JM8K/Q+2hT
rDQvrXKdMyWxo5OhSd1f1W6SRgZp8hyxEhtsAEX4KTINYasNfwtaio1yI91ikRZWC5Q0utyCYzZI
9HkiCxlqrmFtLL4QHcrZa2QsAXAlcnt4RxwyZLgZNR/9hev3VCuOM9o4PR+/Bvj4+XbeVM580Mx3
SfRJTNmg2RinBiftrGY7m8cV813XM10WC3Ubfbf3eN0aJnncIHItfo/CpE80b0Gt7MWa7tYW2ZfK
jGFT5UgYZ8czODc+0+mZGPi4YKs9TMDtIIXJZnyR+pnbZs6woMfQRwrvwC85d5Nl783Eai3vQIAu
RzB98GVt73fKZ8uYhf4dyfGtNR+fHro3Qb8X3IzDgiuYvnl6SO92qYwZgjiBahwm9iCDHmXM/D8F
0jJGEr6L+Ca8/2y9poBMBFfRZ78IPxCRdPLBfVQoum+W6/beb7OX+p8nbVYFgAQFm6nJXFa3xfbr
/JklKY0wIKL+9IaJorBqpdxPCipT7SwM4nzMdQG7fbiRE3DSqWpNPGHibfjmH4PUBh7/br5I2mrx
4XrkrgTFJRPSF8TSQZKRMMqm0X8IyEMdt+TPlIFYp8zAJU1hZ3CwqZMkzqgZX5Qk9kOv4dkPtxsD
ADie54K6tKboPZFOizZBLZ/YKpEY4Z5TcFFU3Gaj1UR/d9t12KC4PLFwN/ZcjXdQTuF5CK6hw/4E
4q/6tFLtb/LeiBzC3zEiBt/WYdFzfc+YSZHemmQ4RZU61txU8m50sljmiSg+fmvfS2KJsEKkFXxG
onPrOAnmqRQnOfna1+Y451QE52nc/e9CTT7eaBAmb+Mzi9WviqJ7NbtxrrNnKfAEA5mB5O/fx/sI
xyYjCmRfT4FdlGbMHgGMdrCHCGaVqjxly9MnQ4On1YUKA3NpeWTaM2F96br2Z9bIINNEIBbxBj37
r3i6OLqXyF9PKQfJkPVXFuoutHrsP5cJnC4XJ+T/gBfC/DD8VVxwhxKnlDtnZMRnf7YyDEGK7lUn
XJIc+DgUiM3NpoBtsDpuMK+/qN/HSkKs0FoEODn9nb43OWR6bhiwZHFt+2/27M9XgA2nyWplHPkf
kNufXIO9vHsCqfKg7CXpmCfwE47EEUvz5MPmeysjnPnjmdotiSrpJ0QnsenqgPtrmhN4u6le3S2Q
nvDnsqpHaFntyFq8sZX8iSThO+e3rJh4HSUg65DGXy2qI7I3Gklyvt+mzj2ScNjJN1U8REkroNh4
aNWx/ItzvytBQ4W/fMRhXFxyH+r+SxQHFv78i8ZUwQerSEVpGsUmeollu4EWSpuqt31X9csLVgFV
nv6rMruhUdC2g8wfiXUBIlu7RDRP1FUPwxVaCebpcpb/Eed/v0q31Stb+z18hHw3DmspY5zMEls/
gAryaFBz9X9+49pT+kSKDr4BMwtQ2NDoNFWrMGJEKtXapTy1lp2fQDQzK76nyg7xg6xc5497WwJz
Qt8bM+smFVd2ZMz6Xr40SSoX+UTsYfnW3RrHuuj5JgaoETLzodHLPxeZhzjGGF7IH6sPBpCmdy3M
OAHV6YnUDOswoFagxG+4rWoG0gWz3yK/m7Zb/8HINDJv6BIZi0e7gHwnB3KEuaK/oJD4R99TMp1O
3v/h53YV7rnZrJYOyl6G3FLafOBrdLNh0vbbsg/FS26+QOmcbnMvwYQtzrRS6EruwikSZH0pU2Vs
TkZ6FokkzwuVoBTCVwBKREyhRkPINzznOwjZZAGcThcsgWGFkJe6AMi8Sh8jpAvj7Qc1kuR13t7u
s2S2Vd/sAccgBtCqFbbRJ8JxNfQScxtp28GzZ4QUAGD3ZmhVn6/zIrsuwTUo9IShOil1Mj5Vyyj5
xd/i9b3ueXPUF95GxCVX+n1YJhM3PJoZUcXMPLlf3MQRHDjlu7C9qg0m7UO8K2QZVSNbcfT21foC
BlHehmi7bHOwo3tBTOkIub4/KPo/3jw+L2UrZmCtoM/NwUgYJAU9UtpNioxlUwqfFdLSQC1R+EVD
w9+48TyhgBcNIDxe9HbqG0afG4wpqFn8ppXVYO+wVw9Kp5qKoSozimyyFnLzY2Gs+eUII8zjSfqM
Z77tj7o6e91xW3R3Y3n5hoyrjZnRROgmOIVCaUYOdjVSbquXT+Ge7U9XZBhyoTqoaW4X0WaybGjM
57CrIM0BB7mqzJ0OQcMUJ/7xMzfvk+ggOJci4JhZIJ+IVYGbLneoaSo9L5qKglg/22D2x2GlU7Gy
rV3FJegLyPN2jybEppXu3AQ/ikYLP/H25DUEZJhGeqcHdXj974TcLl+Jr3/ncwEBpFC2UyjcOKZ6
jg5nxLwDrsFjMkcHp1F4q9zIqlKjxsA/+l8G9EGpmGWG/vDKn5W+ZuwNyLJTqijdouNB/H1tLpQe
XdrA/indrmwUJF4DJKQBpd4AytKRElCkcycSctlHBWie5wKCegvyc4BReB1PxOla6g4sxK6JeoyF
0vNUnZ+KRTVUsiUfW/bg0TZLkNdFN9zfTt7ryKzNjkpx4sN5GUlmoCr3mLLsdZoQrIUdksmSVmWy
bZSSZBTC3zjitBeVfAXeptnKL3oMm8ARKyMdddjBB4t0Ra8pknVJfEud55xInX01ca5hTJskePGW
lGfuFmzTNF/Zc4cqgLaffTajKM+aWIJWYPeur6by8HqiQg22Zjf3UxSJ3PZIksChW2n1cmlAeyB6
CaD6uRYQrEpOjAU6bMxdXEWjaXCuw7APx9j0UAVyipuaBA8+PAjRMoHeiDw5szTLltCPkZar8ck2
qIzEr3hz1f229DRxAeuIswuLPJn0L7rgOyPrBr4UZlGmygvCA68ghtpducmal61J0AukoLF8z9MB
QctdTUQyafNwmwCjNBN95PW9Fv/tGz9nIDoMGnS9LjqYQyWouvV9if9H9pcAxZ+4yKY0onGHYFGc
emfMmgs5m0vW2MngTJvUWJYjwgIpjyvJT+D8GrshxTO7AqWVnyyiPq05Sp7Je6JDrGSEKgA6XreG
NGbr0I7LcNoE2/FgvCUdsoLIXkIkt2ZiRtCbTyeZTotuDALBi6CBb7Yhfy2hNcAQjxkrOYhtEPTW
8hZ79KQZOB8s1kz8fjUWbPvTPc4W5+UrYeEnA9BK+cpEugRvZayYFDfjZKsU/ZeGm6dilx9sTMdd
1VlirMmbCrskSwj3nDVlMOwyB+0d2neIyv1f5O1e+jx179jns9gg3Yrtso6yqSOfaC40eaPBCQGO
bN79XBbk6FPF8+wfbUbG3auw1leVHii/FWz/nljqR4ibq8AN3bmrdxVzc9650ArvLuLD0lwhC+p3
vuGnzqTV22aiEEFy4tmMNHQTqo7dqZMJC9e3RbFgWlg1bLWjoMceGKA4O44Pk/VBxVOy6tjenbT0
s74AF5avbCI6Ag1mooU8MW0LxgfP2o/gXJDD+hHfVZ2jho/+QFljTMwy+a5HT1+Qr93OQJZeL8Ah
yv1nyTKvZX2TGhkhMa9pjY92P+/ff3mtx79Lr+HCmD+3Vo2q2cOTXnZb+JeeCWVzmv7bsYFbEjMh
0lAiMXxMHjtmG/K0vwEFy4AXcGKROG8AewTR5dCb1GY0miNOoz0ivjHW98Tk67YtQlyP0iqQ8y6m
zqpLTYf3VOaXTkW9scfKmg9cX+9ytEqNumB5rXagyG85iPYUMKg6O0iFJwcf14XqFY1434lG6Gx1
mouaIcrSsd+08yipRaIaLHTXe9zKrcuHG6WQGzybB5WIg9z+cSOY9WrtJyrY8tZef6KMMmv3Ywz6
8gdYETDc5VyCKh4NWXQda1o7kfup+fwlo8NQCgDNHdnvbWhtWJZEM/LT8bMbV+eivmMsHk7sAHaO
2R6V67rEiScMQtUHntsE5moLgOcIoUr/3gF3iyhU+v6k3zXj90Kzv5K2vnHQut2PASYELihHNgxW
HNOiI/J/wJ8sWbjfkO+r19syZ3HLtLmbiXCHhUYD4IstUscB02etPuySA5pSHclrUW5qU8HC2qOL
XpM4iJo0URfHAHYDi2H055stN1Y3w+6SIEdgy3j/9gT5L9z/YSyVlNsFksF8l0W6O/i1wL1dE0oU
17jbXbpvnfDnfJTv4IV24AprAd6KvRbVfE2tkjd9Z61JFPQ0eq3NuwD743VLjVVbhoTXE8MCTF6j
a1kt+jUZdjROXhCVvwmpuJtNAWsZJmBoVMPid+F55UijtiuUWKGyyFIPPC2wpQrqaMgUflYhZEJv
12E1VLdsl6egsvfpy5zpYeOFDS+mkdbhYutRSe7zjcnzWdDwsVukA9W/rlZfpXJbIQ4ZAzMRjrEc
ZjDTlvztvm2dip0M9PJpZGsiIurBzHyoprGot5WhqLunkzNCF3hJpiYCcaUvp+uctAA+WNMMBlAT
opqtA9/K9ODo0YM2VmRRWpbykldb0JFajbQ2Oo19vBlxt7Ux58yUTXRPJ50ts68yo7xC17P3fjAq
WOByRZMbEs2ubg7qkZj9bLjhGEFg2+KPA/eik9Qk6K3Na25nO8S2jC5rRqLyMPTE9f2S1vjRuqQ1
tSDXC2rxQm6zBB5TGO1cCsdrY37EVsgaazfephgS66GP9QgiNU2YDJm4ScojY+K/tn5moQIKkTQ+
9mlaKkk7pko/PhtUEAguVtU4F7eZzvbHNBvUjHXn5NILOXePDEWlKypVY9+wYcmO1pXzd+LKyvgI
RiyVDTbO0sVQX0h0RQvSd53CRCtIqg486Pzo9bGJ0lk5ikec2g044DF6ZFc4oNThPwq2ofD4NXC1
tbm51E+bwEvRuKXKUhT5UgYdRXrTrKF5Ww/Wvi06nLwkkUKg9h1LxwQCUeoKIGwIlKcJBbdALdWg
SalyD7/kgT0YkylseFx2+0I05Kjk59pdEBiTmNHgyAfihpfHiNKvsatXa9bLm7+9kA9TNVKRkVws
+JoJ2XTl/+3OGHCFAZGGo2JzKuOKf88TFxnxGiWOU6fhmzwBAwjnuyA6jaF2JqtdZPfJBXdO2j2c
8FreKqLlgZ5b9WIYHXk6wdKrVgn1S+eVLwllw0YUtnEafsr5nMNtbbD8N8AfRwjv/Uq0Emz0b504
UDBVjWbh+9WNNp0yrHxFwgj6tk3oLECMwOV7bcsISsNTCeUfCKxWpldUzpgvHrFf5jHmKrkD88Ab
amb/fdk1h0W3l+20lxN0gAF05uKAi9ESwsPYfHjqSMNdNkR6DpzO1IkC9vxEtrd+e2//khVZw3fG
KqgL7Gluw95RW5VssK1MXCL6V+gTqqr1xzqWOtT7sikPXvuASMMCn+dmVe/C/w70GYz/FPiOR900
8rNRbMTtMCFsrGzzM1SK8AqTNNYRG1wcz+hAXErnTgiCQEkxcc8BXtUu82g/GV8/Y5HSWtq2J+OD
tHDfsfgGxCylWcyS2zOZ3xu1EirdCKcXu62pKt/obMZljq7YnqcEa88TDibBKUzjKDLHsyXk8csl
GOM8aM+WEZYs5gqK7mAexF2BV8NUQ+shzwsOQn9WhQOow1pc/V3ykqWJkiCJsbkKbjFmO7o8RxUs
ObZWnc0NOjchqXwR1TlsYSo8WnSDBJlmGu/fT5oHm82oXsuyEqkJveXPWwOGquKPdnygrHf1wD9r
LSnZVsTB6L2O6QzfoZ/QUMhC9tws8WRZwNEkU1pVZrfrDX2x8ekzPv0jF9ueKfXELnTtHmFuHDqc
DNVH3TSPLcI8qxjl7ANIA3UGIK+M4KQ7BdkyIYJyymLtOyEjXifSh7ZbHzTIIBP5+db66ztkLgpx
GBQUedQ0UTrZXXny8QDH5iFUR4+/tztAV2YZypotUL/kYqiAVnWQxm0DevLUdxXE+f4ClVUvWBKX
sKEKSlL1umpV6DrC0E/0ooA7BI4jk7/hBcZofTtB9ayFobGl/9/r0Bcwha+JYiDEdqr4qR5FeN/p
04f6Suji+VQvpd2qDxZliDuYtMcETrU/woGSl6doZ34oSXWZlY8U3bC6lPlmNBCsfR7P4YgAbM4I
4FZfTyJ0TccDmVjQDvzW8ZkLcWN5qnNRILoF+unn6Ye7vDxEVmwpiA4wvB7GnvdJyX7IZ1Uq/RbS
7mzy0lcnFXKPmMy83ZtMgHJCzGu7rE3Wgya392f41G0S54SSXyOPfMZIe+pwjrw0tQWAwQusMgMC
01RrZ2CpAbgYOLkrLwNLBJQdUE5upOEAXOjU8NwGTCRyAcpoiZxLxZdi8d5wMyUWjmimkbx2ETFt
Wj5FTEYYCzPWb9MX9v4dlqH+QXgk+OdyLjrdUYRc3uyw3/y+pjICyHWpuBkL3pw3QUWWGgnZcqVu
qsQ1SrVaRHaZ/k6G/oJQOqkNsY/1GLwxsNnJxUIshb4shnGrKFfuxZ0uSycVVrvN9+8AIpqDR8eF
CjJWcjey/M7be3ypQH48bxwEgHRqefQfDQgF9Btmyxp/3M6e1mr+dxoSsnEH3R859+gXoSdbB6On
jAXk3REBto2hWMViM0JnCYnnryjEbfWlZjM1cPkqwa7OyXKiMD9mtBhuQCy9rVdf3UCT0sZRvVgw
3JIk9ugcSK8nkTjijht9Pd1ZRzQH5Oj0XpsQLdrdy+DoXRrvyuW8O4Hk6J+LJP93ioJuQqf4lS0Z
o5/RzECClHqQqKmopVFrr2hZNTg1BUxnuXsZK2Z4QvOrRYOLMqYHIMQgK7+4l1DGteneken5N3w7
q/3i4AVlkWm3BoD33c2ct54wUcONPG8gwjKfS/wKS4QAtRzKPTtn3kChvUOdKWa3T07l0B8EX6XP
RfBGXcUmKBYv/reSQRiM/M7ULXFOG7xEKuoQg3LHTZsRtszXgpq25u/C1O1bxZ9JHFQ5Y5SG1VnH
oqfFW+EZz/ejK9Vd6umaryNxlFJC1t2FN5iPJmSyoEA5T3Ux+LJLw1WH1p6qpLeSGwnUhkncvN3o
STPYOJwPGejonf+teKem1BqTz8urmOT6+gkGr5amgXkP1SW8QyJ/XySUmwcmuFGAqYqLh1RetrPV
ELb4YVXQrscj2lUF9BUEbwSHaEQONr6DwRGiIjOcPgz6iWxsOtY9X5jzKTqCgTbcyOWmju8MXGLk
URSk38dvosVA4qYEbp15N5NWCp7kewiYP1IhztasPyz3l7WuhJWaNv0WF+PS2H2a9w0PBShUVa4w
jcQX+Eio2m2lkDrQb+CRIm9/nz1qz0269ZYMweIEh8RA2b+39QB8JSDlinBWL/DDpEWJfnkuj1QM
ylcSuOkMPzVklLDHqg26o8z82KsOQ9hm3U13FCXWbULnPHyijIU2O8iZrsr++C0rC3NvpVgTiVMX
wr6fmcYAL0G3Oxf1CninhbfcI4xlq1IkaYExbAN6pV9eT13nUCS9qTe+8DP93tAfLZ/rnTUsR/RW
8kdwNWeKRTeRCw7hpWrmpUpsifMYqhfT/jPwjYkbMymLTKqB1tILqLAWgVAxVp7zyc0/2iAxkGd7
f5v6VemEcG8zCP8De66/PhqmcgOJ5mYH+eXwvcIoK6VHrPRgugoIr370XUUaiLNy/Ae63BnqwVGf
R2STyXi3I+vW1jU89m/z6IOtmuvyjpOlZFQ2e9pe9q/KxtqQ2QvI0WQikB8P0wCT/LcqiXRv3cNG
T4WnhvYiok+B+e9ei39tSz26xV+jLU0R+UAt/eZ+DlFnYvefG/Tyr29NF358kN4+mOxvALLfltUs
hjt4z2z24wUSTiUpmkSV/ykhsI44KMcEVMlxj3Y6au1rKdSQ1uEjrw3gIDRoLCN/zi26hOoIgQkN
1VFw2svlGQnV5bwjBF8XMvr2J3zjweUsWBxE7aj1OeosglDAjeLellM94LscnfL9Il5yPWQHNaBI
NLaj8hnFMRDoXCS4qThr5AVp9RwMgMjjxLdBeBmDnq8upgUZJUak1HnA5lMR2JqtSw52+hS44jsd
TY9mbXrbDfPu4tGNySr1v93soX9nEUeyFma6UeN/heiEcYhVQdRs9Ykcs0spyQ2TUIs+XV7YN4Bl
p8OtvvyCuvM2XQ8TF+SFF178Tax+TEeHfvnRmLaSh7QkkcKte4xv9zLIHYEbr6f4jRd1Da8122zl
QvWwl0/xLizMAwqvkQD4+wMmUoZ/v29ZdT6rv3DmewNXt3AoVI4LshbYJOMv9od/P21RXzt2LdmX
HiwfyidfbGWU7yUa3IPfainVaBJqxe1qk25w1djXyrH1SJjPaRgFwiQyDWe3J9LOb8+uErZm5NkI
9Aj3sjWhkiWXASuU0rRztdzZ9nRqZ+YSeWLGi2/r9LVZU/Wb0LtscMLQO5xbuSmK0hWb7VDEDEUn
JN1BRp6u6XJhaXdBBq5POPhfU2kycfGtEWLd6V7kaKlLvNkTBb7OO4bo5NRzVqyNx7XsuhqI/ypF
T6H8POUymRzlIgHHhCCdEKjILTi6UlY2NB6ewVWS2n34QLhplv2/tsSqOSC2qmu6Af22p9RWbzro
XaLBhiXTTsH3FDM9TURj0MiEVv+IKRE3wZMBH7OQtoLlqSRoGvuGMaRnlJAoQ/JWFCYUh791k2RN
/3vuBDaCTvBl5jffH3lSRQA+Gp51XSB8FDrFo12LNInjjZXW+wQbSv4hnheoe5fbJlrj6VPYyCw/
AIfIytFEadoyGrNOPsFyPuSk2+3aHvwJW5M6yeb25dhbtSW7aUZKK9hjietExiQJfl8LJQSFt+ly
UayG4tXWqHxEgFzvHjQnX+QyprJ0A82ntZa6eRYhUqk6TeDKuXsvitHfSzNRGg1yrFPvaqRSJl9B
1yXLEQ7ilsXH4L3VZ0bhvhRVNW/urXsvUBGv3WMpCedg1/S5JYOizwuhzxsJ1NFAhJ2FkQlJqmef
MZvXzeDXevCOsAMiCK6LOQ+m8fqlzh/hHGbSomOWeHCCbHu7HNKtamL427oLb3MK65ZVJ7kc8flZ
fgbOAiYgbSpcVtNROqAsEPciG4wO0PaxLl5IYJu9O6w25xZFIJps/n1eZgZCuMJwSg+MpGCdoSUz
Cfwm0DXAJFfAwwXZB/in+wl40ns2lEJUECRsgYo2/nCO76XyRO30vLPtPt65Lmft9DnN2aH+u4ur
DlghssioqqRJawfovihY6Vaw0oAblX5smC3/ow70mCcGnvF0M0BJb6klvMkUKdiHm2Wv9zcMmjho
/YcgnIjKvUVYYBoUAqgNFA5sPDmG+klJd4wNBnaQx+JxmCKkSxVPjKsVKfhemWW74SgM7FJUNLfw
/dPpH4dReJAhG20cn5zYFSXecoBsnvvBMevA6PGqXboiZo0iwGFoJwrpScEdNvM+Kze5rkkqlGDV
fSY8RSewqI49vVUw3MEGAolw3AFdiPaQC1sfGuvWzjbr4ym7YBQS94YhODAYwMucMvkV6rJxoDEJ
C+sXRMOUtmAvXOXIJduM4CBzaC9z6muqpBCs+WLYXn+2wmBQLv3u2XOK4vmErbwLqAPRjxYbibPa
cVQ98WJ9jordvPZyaXReJtf6qQmD8G4aDjMSj1u9XXP/L2EFmQKbxbYlJLdhoGPbq/XME3nxIVUP
2BH7CWno7wLgAA4WKecewwC90YzdLZ2AGcFJUH+zhiGlx7gJxLShOu1Skaf1PXZngTrTGfE/ibgb
4h0g5BLxzeDMI9j56CHrvihAb9JS9a3G7mYLmBZuBjJOCTYz9rb69kBLaF64hyyfs5Fq9vZWSLzW
/OCflNBE36ydAotn5hyB63gOagOCaJic+fIBq8sOCJehqP3veIhQ9UJyc2XD4uUfC1qMiAX2Ip/b
lH5w8iEFurNJRIXeCphCPcqS9H/UyiMPVi2gg25yOp7rtFn/IIliiJjtfS5H2ix3c9ny7Rtuv4Za
6aZpQo8rP6FxkNWMqv86eScKJm5r+HrK+yQmwfhQQUshhuHqB3RVSyPFeDt7fHJXpXGFIugu49TT
O17Pnv/ncpO2xwFWOgcisCQ1I2N8WV+27yNywRjpo1zybrJrBqisS1/yYGN1GyGE6sbL0AgKFbeJ
epNyyuChE27LG2RRVA+UTK8I6nzJuZR5M2WbbXWWy2Fm3Vn56CvSIIGix7fOK38PChr6bhGweBkj
n8QY6VL7yDCmfUNoPrJrWOltaJSM20QPezX8l5gx73rrVQ1f/asncJc1QMhn0H0Q3cx/zw0JBAXC
XBd7XZ7qrKJk1bRxM0r3Kz3smDeVsTc3Ee8ZCZ7s5Xgs/UPJNYIVvX2oIeIKrmxYZ/LK0Lw+MUtf
e9ReT3KZKrhf8qYy0HrBriPZHvXle/5xUFXw/Rot4+sWsD7bu1xOlTKo8UiVAGdpSy7y0eJWz7DS
2FdC6sevbCzIKjaishFHkgnUVPSVox/EoQX5RKKyFCm+DExBTrP4+i4NnP3fnJXiH/8He/FBF0Ns
tlFUdPbsA1FItyZBXJBgV3o0eV39ReXczgHI2Jr8X9Ro/0GzowFhOvwLO41Til9bgPn6OGgho9h+
R0AtrLN8iztMUby785mcwM+kW7AiZBaaMWpdtwozn+DdzHe4Kee1pVVeN1hOMVT4kRzOydJbfYPz
i1e4dcBKcu5NptOdrm/7rn7EqgkcFyjg/3gQraJNLjb1XW4KJxyD6wLD0Y/cAEG7bn7h0nIzHibN
7j3G8fJJpG6AGdwei/alih2eFfZFgw7clOV+txzLiUZNGyFUcj/WmyVd5EotIvvKFUgyOL5TdQno
At8SK6I4urwOtPw+dHMXwO1ewpWYzrh0nrEHAV5fy1v7wfYy6caX4RdAAjWrvo3nn8UFeZP1+kx9
+9JQ/JsnHnO1vd4ClUUrpI6ZwuXADseX21+wo8bUHK91C6koMXLPBckWzWetu+4L+COB49UbNxXI
KW7CkKSxn3KFC3lsD/8UK+bKQM1OwRmzl0L9043Ph93siDKuuWHVoWohe64bZ/9ESl1yPn6FJCeF
9al1AbHCnLrZ+aN2ygsj7Xc1oYIfJJxt63kmEFR3pEqEYq3sm99tmG+CEiPfSqs0oKf9NNOqNcOb
6yoQ5C8fAEsmuXa8chPGECJoc5WMpPJTWeqgrlP/6c5DYBGJVLvYXRd/47STf+0ZW28R/P69dFyu
ZiSfzV410QbXnu4f+3e7QH7qCWd9s3Zpl20/kpcoXiD65cq6a7pVo27n2DoECT9TH8/07VmRrt7J
8+CWKupQ3qKtDNiGpLD6rSDtxRE/n2PbYwakDFIv36YifqsVL9abecK8HePomlOFZvc7nYwPDu9s
OzSl7RMxPrvujWzQZMPhv+BCEMl9joPL0Z0Sukszs8vvA84Oxi76EKi47HValoXywMXsva7DzHlG
b7hbUv2BRisDdAw/2jREMGb5E+dLgK7WiDuVhbtFqNUmCYAB6HjkS6UTxdrobj6/NHzFhCekV64e
2p6QFD7RRmZ1H5N8ROQbNSUt6SKuBs7wphSE/zXoKtSWNmPItQFfoc9DDiP0JBdbLVFUxV3SvZE/
rLXhRYp75i0lylxB9E90a4XpMJg0rvVzAGPkUkdj4EXY00mM2erqcHM2cmWNF6/XMHlF12z/c51j
u7AiUoSPCAWHgNqHm6wQWmxesH4wmXlifaFklJYYm52zj6H+d908Ofs5cB+Po82+bu6Vq7aRdzBW
0RUA+J1rTI0a098zbkRKISOO/Nho5s3yJEUSbZkJkwUX0rnaN81Mq/CB7HeOPwkL9Rfm2kQRKl2G
H7OISY2WvLraigLu3vUs
`pragma protect end_protected
