// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NDtQUKVw8ZP5rEJ6K3rCbH463oDicqAr6Cgz5ek0FUXAEsDZ+Dk3SYOCpWtsenSz
+fs5knFjyvwW9o3JJCHdMJIjD+Fhmz3wyAcAWO7jeSlGeqomFWIW5Ws2+InjcyFo
9eWDaObW7Tw/4dhGufOw+KqlWYvTNmLWuhRpdTkrH3I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58352)
JRJIu/6x/DXNfZJKjg+1vwbhZRlQ4rsMnKDGcYHaWHEV4V067ZT8h27ddiLGAxy8
xPdOS/rMpc1idSjYO1a3bOvIPuihZ7mSF0U0GiQoNpsJzpQnods6904jue7/RcDy
bl/el6RPuVhdkIWJzkjxEfmS53hQY57e3Voz+0VWN8V3lohM0b1lpx0f8GKj+sc1
e6+OAzI0c2tlxKuArphPC/Ct+F9tecvNhk0lkMcxs9A4eXL7AHN3NeCqrxaOra1G
oxUoV0lX/2VQOaAtJoDC2y/zs3NBwa0YwhBV3iQc+/bxpxNZQ52hhCAP81Pe9QH9
myVxAdhQ4h+3d2ZU24MJ6jWEFige2uRWzrk3hneSBw7dbNoHWdcJogv4Fayj6I9m
nIsAWfVAkdEgZoCv8czVF26hCw2eBpfgEmrAl0GM8i5UQRikNfaK12E8kvppKqx3
WKAm5O+7jOKFG/A41TqVYBnXT2NsbVKuf2llcqiJOht6+7O766XX1xyNgv9UCRTK
tzcx0jmHWGksyCPgguEDcMgh7QjjtWJy8Zhz2NjmtXMcNL73n34xTgmjY9mCsMTX
6EoWPnY8bIfZqH1SxP5mgTWUWct0mm7yDXD6oDEfO4uEKpH19L1qiBMpXL5s9fWp
/MgYRV1L7sdeNm2GnfIEnGz2RoeoSD4WDoDrhB8Hs7VxJJOLC02Lyo8V6twASnxR
M7N/7uklsg0AGE95WMgASDoH5IOmf/dcZomPGXVLQ7oFt8ICEEmxn5wTvBwUiCFB
jxYhrFAyNqsQKNwGZLzvZpUOkr3mZDbrFyVD2lnZLtJgsJPkxlPuJI0cyd+21IyY
O5zLgTYvJjP9XNuLnD0b5qMUACs2cpNXZeZn3Nh0ljWds0Y5BWUEjUomaTyRj4M1
gROigvHw8fG0xGaVeO88FdRGotKLq49z58HQImiWv/gj7wGQ1WY/LVmZCPFAMfM0
SIE4AWeNOiTGPMSHATow1344wvjh3xbEecvGp+nab9wAKU8hkJUdBn5jQkWwVz0D
C9W7uFfHWRNFAs3vlbtyjIg3VDprmhs2jVnKksmL8T+AGFcYcFQFFmqcYozVTzdl
miGHdg5gqZ/8n7nP9ovshdfxXG/y7UEBN6p/j2TJI/bewa5xZBja3L0/pEb8hod7
T+3lcz8WJ9/UYgE3dGZmox19+yylwLaHc7G1zbj0H0lJNpgjEheCytavf3/elhHD
ONL85OClsASLnxAPKBexdwsqyJ+7ZtTtfFb60dLSpt4gwKPz5LoYCDuiAi8mxYTm
+aSBalnkYLv+zByMAEzve0yNvogKh2kvfedYjLhfAhLSvBOhktGkMxBKzxjS3iNR
5fLlUdekCxEh8rjiSNI9ZoWkOU2d7Db3ir3HFV/CJ0cFboFf92UomiKJ2ASa3Eun
hXC5UCMQWM4gA3sQaAEoQ6aPtyon56wYQ4YJPQXrhkF0FLpj7Oz2BmKb1TaGgEJt
M2zByHFP7a+DgxALmsTJJRzdCoVB+H06V9RwlSzzLUVg393VPODrkgwA0EN2HiCN
LNztPqpN5YjR6PAEEqbWK+yBU+sJEG8EYDzjUdmOtUdQtVKyXrfJGFlgoP+J+J6/
z2rQKlUCvdNrPnOaiqAkp0Pt44B9RmyZrCYVpIFxEsnB9qaq0V9Au9sl9/Nmd9pg
0y9dmYOikoBlNOPYFVtzRfa+PZRf/wiDSWQdTAGkjYc+S12rhzQhtQiFJ5tpzjFd
eHJBb0DpeC+dXC7KLO62hRKV4+C7+LYsQcbSe1A8XJmGxcEapq1AySYRHt7Lkzob
XyJYUK5GZReM5IQkV0JvKb2tlqwix5g20r2mOnDXA6QeJxfiMZXx4euxyhsuWqRZ
DX8AI0LKCOnpaL1+JoUvB+ouMyO1oK8sHMX6fkEaYW/SYA3SI7S6P61CQM6gpw5z
gvY4d9OvCpPWbV9170B/gaes3GV+ZcHwo/WgSblYgw6JEext2z2UXo89AjpShyQB
ks8PtzfmfrsltIjuOcGZvHhofKyHW2RHSVA2arCMTXPBQ9VKzRnkzq1DntBH3KZ5
yZlrv5TsHm35oa1qsYj2gwTblVkcRXzWWC5dpfWAlbaL5c+nkORkZGRDH6qh5zOJ
UG4XuaWeCUXz/l+93LAq7JwwmULHvaVMWWFmiMsLnPjH92/raN/DuNaE92eEiGhf
UYM4cj4Wyc9+izrX5Sp9nGKJffp4Ven2YT5GjdzKq241KHFTenhHH9LA4ozXdnaE
rRPbzT5STbTijyHNVfi07zsMfOEtm4RYgdXOfme0IJdhVv6X0UMTVancwLKkkxqE
qm6PvfLrMcu/VlbsbkUDZ+hrjVnzporEUH31fJk+QBx9ntoUcFGARKZR/TkGDPf/
86cxaFretx4lkg45F2BQ9okjqYtxgWhkHex7B3npIGQz3Aih5dif+Qv/r68sDSDr
WXWWU1o4UDM2PWfcr5+xde1yIf/Jys+ep4GbVghScZTPhnObHd66DExpOyVkQ+Lk
hwibEz6rUOwqbubYAnigrQX0sqtPtme2/GemcUJsvntaFQh9qEwLjcIEJo9VOsIV
mGgGLpriX6QO8P70cx4KYXvRt6VSI58LxMP+cFlZV5FAkchR8CTYLasZxoSPqelN
sq8iPhILo55Vz5OlOxI+V9+hh5hSG9RXCx7Gs5cacjORWcd4XegDaq1PfzseI5k/
OSUt5RTlTCghbUFt+V4f9HYq1zSPPZaXPHSJaKFKcSfumZx7FZ2F56ErUm/zCwvU
MMFufTzgE1JlOFPPzWulfyE+kRRoiRrwLPf2ulxcSI6jV9A/i2FB0DRcSNBQgLcY
1xxapgruBn9u4LRN57Lwvke/tCl5gn8CSXnAtclyHk94VJconc0VTjO3Isc/7baU
33UtXMP1odC7hlGW0BhxCtGKz2QOYneM+WaRE7RyTFaaD7hyIixs0N6pUjQdQ7LW
nWGTt8NIOq0cgAlfkXC0ENxf6uwxxrAafQuyyXB/pUn53Qxp87XG1Z/OoZs6QiNC
3wsyObHXULJ0UGLFTNq3JhrXboQFUIkN7cDKImqkdYBH7XI6JTD1/vJlnKZjePsq
l593Ji8QmERSHasjO8HJuCoOvB3LH2UodntDzgZbWLzFJgavBBNccATavOwp1Fc9
JidSnpE8mlR2Mdpk43gGLujhRIuv7xMrg785yHX0SlDJ50F9/rtrGiSYtEH+9O1S
baA/tO6wcs4u62XldYk0YujVC0kcbr8ToQi1NUBWy/qC4tjeghhaOYeTJbfc38Gh
nilsLnch+0hOQM85vl656yih/++nOtmiYUgjmzw5UicXrmlAJMaayCwXtoo/et0w
+VDfPiz5fJ6A6PbUpl5Ns3QDPAjYDIlLZUXRiTT7odmV98AqBg3OIYX0tlePoM7n
+M1SDEpu4sxiRlzqBVEAdwwMujxqcCiw6fwuqCIN1zWdpmkCI2jF1Bjye0jHLLHJ
kU05WkjXrrbpbjf6XNda8lC2hBl5aA6X5uKqBEVtSRey41HBzzizYsFPGW/qHG7I
6UN1PkuntIeSde8DTr3vL3QDVFOZ/zW4Tx41jMVeSZG93wfzc7EThO+LAUmp7Z6B
IOXMJUrySKnjbpwFQipknK2oIYdIl3i0KTRDvp3DLvdBJorQDWH99Hx1lfu95Vpr
K+FoRAg+TtysVz/kTN/e7lKtdqJReli9VocQ9Smy4B/DFefFM1iDw/EWkmd7Mttb
JDHJlVcEyN3ieUMUVR8P6yFAvM852eHEYK7MtqORxhmFEHNEUmiCu9al7Sm15Cw+
v0LqiUc1OT2zjhsOzvAlSoL0ZrN1XK6WYOtNbUsQbHNiuvRnrcAuhSU6sljVORqy
lDxHzvoTLpSnEwrH0vDjlGKFKks6vp0IJmXx2PmSX06cL66GTsxnP1YItnyYbgJd
dZ9cP4mjozYT0QdwBoLUvl2ZQJ3B6wZusI25nOHPmcA4wRxh8yu5eMPV0hYLtL53
GYW0ENho0ovNgxYACrPBVzVmC/3IfnJmeE0++ObqSy+DJtcwAj6oUVj+NJpauAo3
G87jhdsdMn41E/ly3KB/88wwWH6OSogk+elj2H53pyrX+E0Mg8L22UORsfaMV/w0
rwp2i80rs1m3/yT5ueRBFDKAgJGAB7YFSYezB3NGuRwqaShx6MxP0RxSXIQ8LDtq
W+bhhpXeIw3VZMVmoC+ywB7saxagKCvHZw4ub6dGQUOnS31z6qexaeF2PaGwZoxP
Q4d9yOw98g9c+MK2N3zD1SVMTG/KTnYetFq1EGHTtqv4jR9xGWjhkeiN+AShJlrE
APdG44i5ZSQWrUGmQTaUMR6cG9VozcGloG6ql3LbF2WX7lEGOKrqGYfLf8/qJ2gw
cVPC/+ozWpkAoyWoY1ZXtuZAsYSZNBu1kXCQJPchroWrQJ0gH0dGmrNopZLzRFof
zzyiLe3vH2T49yIIPGVHP1+Wh3gDFNO2fOeWf4FoB2SEVQ+ino1h3s2vPqm2Ejl4
IU7D7ThXj+lYWVQMA+jARfaKM0jJ7PtV4xPRFHdHE5rRKXW/g0jaeMIMR8r8OhYK
mBcv444BYfVHfhEeiH950ZM6qrtAgt9f9T0uQge7mjVdYeSGKwgPBcYwExR6VeM7
2jB/gNwrdNvi4aaW32XO5taytmrhBQi5ymC1s0zWUh8KmmPOGGgvGZ6ORE/qwR7T
nqm5VPR9iu0/OPMZZIRIh3LZPo07ewENrJYc7qIdJHIOo2C3JDqsSueUjlxi+cum
MuahjnKvVVfIEc7Y815D5Y+DzjJ5NBirf4jITCUj+lB9xoDllDex2twRr24qwP09
TnouWqkUNTIR73wZapF4eURCNPRpaxQ4Jrl0Bd4r7eL+/0cmoLv6Jm5Gq5Ed8QW6
OKc7O/xI0M8mu23U+JhpJwEGihMhah8S1/fb3gyPCi6Su/KJOsCYOGN6EiSH1TWO
2faeKcu32HZbI03hmqm5/JnTnD0QvQ5ARbpl36zaxXVKt89aMz8OXVLGtipcaD8+
gQUotcyReM9hPfBz6cgxXiSrHtKGFym7zyAOqmWPBsAu7gloU3xq5O/7Qz8sYcWZ
TfKMiMvvsStVqPt508tYymnN8FIc4S9YHSpQIuax4ckwSJ1iSj/IGpDQ7KkyWLlL
+6RRLiGFltD24TRCnb1+Y+3v7hOVFB5Kh6o6i+7TisHU14unKsExi8NwcdnEQHJO
9Eb5xdd5/RXR+sIU35bgiYui8WmgGtRogpfG+itanR5SqMxe5N0pZMm/b3KcV1Mj
mzHoJ22ytGZdhGkd/4uXmnMVI4ysPfy8nJjMH7CMKPUKm8TaRUEKoA2LDz2IQr3z
Jf9TLfCwQ1LN9OqR5Rt6hVsxEvwlg/F1vkRDJdPrnZgNe+uDwk81QkuAYPUYdeyg
vKHDJKPKh43MtW4BuZlXqRxnwGS91EFE2cNCRqsxlzQ0rB1nz1ChpYRKw3OqNAMv
Cjg1nQm2/ccQOTToTpeWbW1NwVCCWYWC94NdScKrypxAiaLAACy3uRKB2Vvl02kC
t7MFCRMrgoGz0+NdQ3mkMrY8YCDzGe0NkTmYBgyKN362SdpySVEIBf+ZZgsZ4zuW
sjsrqWWWNV6Xgt/isM6U8RKoLaEfQ8aRjEEtJo7SmiMXsycUwvvYQaDnS6PkNxMT
gC+lvjoibihFJlMKSDdebwDtr+N2aaoopO6RhdnXHHB+JxE5CL0Hpn+TOrwhGwTC
smoCyr9qp1EcaRE+GTTAn0guRfkhMBvWQwPnw+tBRHcMCUPe95iI59Xpzl7qMw8B
jqM3ciOyEmLZ70viqbgHkqylKFkfaFTWzClp6yPLD+M7x6byryPdbLT6M4iqYEGx
dep/EJVZ962A63UaF0yecekcyQMdyl4i8jy6LqXghu84lJ0RR73gAbwkE1hVPSVo
khna9XatcxBl8s8IDJLdHAC84h+k0BxUN7ZbQG4KIGKBk3ZnmUBdlG6O9fl9jc0P
5ck3dveD9xdhai1zUu13hZZH3UkRisd3s3AKll6gWSlgrpfUyZlchM/B59pwbRtb
VabHvfwQvP5XE8lRFGhIe+ozPhV1xeP50hWj0T1jMhwq2WcearM7aW/4UYnWlzNN
ecSh+Ngk5kexBuPTFMmuAxfLveq6BR5FQ5RNfz32Z9ykwOYkCPcHxfS9BEAh0t4Z
6AKIBCxviT4M7mUhURRRdIXMAqTbYQT6wIPrySBT4vkc0aTet+ojEObMyizx+nxa
J/WS7MsENjCAH3HnM0QJ15kNlfk4YilJjZUP8q3L9vXUb13JvVIROfZLQDMUoZ7K
XVLRHwYHpvsbj9tzKpfXsTdwKi/eZqFjmNennJr07jA9tsINRtGqrvM9RHvAg5HY
FlRaLCCjA1A7ph2TlwzHdlbnSUMYE4PNs3m8+je1ijuah1BsK5rc25dEUU15t706
lNMSwEcF5cG/8eL7ijEk5eZTfsF9elBCGSulB76c1TIzeRM1YSlufm5Hm1Xakobe
LRaoqti1qiUOoQh1Yy4FKYDgs8PsNRPGIqHUTC1Iup3ssW++cdfLXaiHrshmCIa5
kHtlJO5fbTupuSkOx7G0zG4quKaqM/uxi8NaS1thsIA2eJUZUBKlWl6jHqnHttts
ZVMFiyMYb+zkhL24jXobSFEuLcC5zj3R3q7YQtaXKBI4xq4XD7yWtcga7qoGhr5s
4xyZN7fWRhTQXGVFBz5jV2Sp9DNoUpXorR8dMXmVcZzotYBlv7CZdEeLo6oItqdB
ngUu7L6JSa8OOJRnrLnQK4xJDs30BmPAJYqYyzO4e6FER5G0w3LiroGmn7bmydBi
sX1etVaOqL7l3sNMKlFnO20GIzq45iYtVeTGhTAEyx3Kf62X8sectBBztd8p4uRu
Kfefp1j9JDU9yuHZJWVZV+qAsSfwkJ/UMvbqipf+FFytvPildfh7OlSfH25MgJi/
uJMnt2wvbw9JJayBESuC0mDGd77LoSqYQQg1iNLG7+qLerLLveLURh9gr39I5xa3
lPjxlsQU9PXM0QAuYk4oAJxMA50SgVveI4FauqjRF/8gDS1dp/MWv4UrGRJ10f85
dwgLswXFE7PLkVuSlFdX2lDzMJEoKCIt9v0/g8UfZ63O3abe5Y6dM0ceRxhxZuIe
lFatT5oanXUMjzlmHcaNYl4Nd+5MIiPZQUi5Jj2lBRqCh9MjiczJkDA2M1a1q7V0
mh0p/U5z5EFuHD81I7ESFId2XrIL8I+6rprO7ZpRS0B139ADhHfqn/mP8wauxfST
vzuKh5Om7/QhmTTv9pzNNkQC5Zd/jzTaVE65mopnJSe4MYI5NC02I22WDk/2eaM1
irH9VbrUso4GUW3fnlgh79sBEeOR+L1W4kueyrBmjDpXVrUJrBWf2hDSmPYuYt3F
4DtzqoLDSIVsuNP99nMwGMi/2U5G/rApbr4A4oQLMIBu5qVM7ha0gjGsFhZKJ0Dk
A+wg1VFupkhQXpWOKbjqqL4vPxTl7xBQN8AlgEbzZpEbwp1FvQ09bFFnFFH4XQW6
aNR56b4J5WjeYgGlwgmnlTIrLesO5Rnp5ZAfJqwDqKwidrjFAOWDmUHc4j6SoIZt
myas5XQLf4YxTcsB/uDvS9UsheVof+be7yr/CkJWiQUtcqSkAofFeaU76CJL6Ct5
8CZKdTpz2ctmED7X3NuDcqUFxLdMLh0c2VdpSIeIyV7dJZTdQMqaCPYcqJZrAcqk
yzW8Xm5cg5exTBP3W2/01nKctzKZVg09sOH/7I5LkZtie9/s1hMq7tX/kEaceJW4
A6Ufqhmq0LIdw4azt9PR0cxtysMqqfSydybCadRBLNeRfPQGJSZMjXi3dr9MSkJE
JtLK3zwEmNhnownUlcdtohfQfIguaGg/uoXOKMXwr7FQ/AcMaygSKOzpnKRjq+vo
Ew6WEkXwrtTR9nVj2fwi+Eb0W89sXusXkE8at5e4msW1E2iPHdm/tLnlW+b78WTE
8Z0KnAJxYTga8Plxe1HYSdTElnMvsXjPW3nnEBmEMxcoo8awCjiil2emm8LbAARx
SeXs0mAowjfMfndgaF3Ze7znHcOKo0b2VmxeAUmasUFBeNRug1u8/yjCrdEYTuP3
DKaPhP+XFdfsft56dBHoIdBLxg0URI5VyOb4C7IVfP9JTFG/atGHzSO9/y68q7IX
YTixYi+IrPS6eugsEOY57n94l4//9HQhSdzEW+vaoes/AN6GAawB7N+D417KBTj8
SUJrdEa5bAIvzqbBiAPH6soX0oaHFB7KUs74lIzZrQz1xcUWvpEK/Gu4HDAcjJ+g
1iNUHewDe5hpBHYcGj4vIsiKrf9RdVzeGOGFmLi8odwytl7MzsszhbXSCa7zT/Xc
fFOlTLC4U4zteaGJJIQk/c4P/noLq60Yqs5EX4+1YY5a2GP2DMb2MvyiGdDyfuXl
fLUtlwQRqj7uLpMLtpJ5Dz/Kmk+q9R5aS8IXgXqqCC5fHEU5IkYl3+sUdgiZJYUb
8t2+v+yc9TJo9/+0VJmkZZnUXzYnzdfX7CVSMeRQBlj2tOT7Qi4P1xOWBFmN8wxO
n2E8unFTP5zNOy3rlp4D1XMxLSNL0Xo3bN9X5Q6IVhstxOpPcraE80AIwZQUms/l
++IFqN3fXgPPwrlg3tyv2ZwUsX2FQpjOhN2ibV1l6TouSeFozX6HZ7airyBZLHC8
oVUFJyrQd3UHPpSPzqFXWgPuhSWaZymuJZGlGxcwhrx/Gwg+QKX3ooPjx+zU6GKs
YQya0J/2inG+2khy97M/llzHxsurDcM8LY/pHUrfXuk7mNxOS76F9jztrwODY2zm
gzLs7YOjfKSaqtN1kqcahU1MW/asF3+VJD8DzykFGE80Ll+3qbuTlQDM+ugSJ4hF
BZ/j9J/3OaBMik6uLH5Gc9q3jjtWrd5Bg8tX3cecY+qFeGpaTFA1Ix/u+KwCIcoN
pTSoK0uk4EQ7Lk+eD/ZL/B0qkzKE1hgpk0nBq+u7QxqeiMg68saqWdLt5rXO85S3
cRViVXBLLUbOIWYOTdivskdga8XiDQ1nxtW+cEmzXd+oPMp0tZOunOVTrYhpSOr3
keGgFsw153C1+cnlLJ3EWua4Nw/4qBpdK/nioscGo9jiVuX+OBfO2f8LRxomK8xB
YrGbb3qCfaV15R2nX/c2XsBoyiOwQHMqHnxMtuKfrUQew4GvzYK20VpntNXwcT+d
VvT7ZlnpdEfgS45qO636srW/yubxS9DsxFeRePRSlDzVv96GYbM5maudbDe/nlZs
Wg77HsnPueKyPx6KFThkKeEm+WS3MaO4jc06FG7iUh/dyU3SdzJ17KOQEWxB4ziO
vXxkz1TjHlKlbBQaLgwQllBLiXcXsYxQbEPQ/U0avJFaLqv3lHyWT2HYqqMbQIb3
cBpbmJ65fmucvyr2HysGA0+XYZ9YzpBFarhmLyW0lcLKHncc//4yEZ0tSf2enAUJ
R3Vu3vqeCQbbxuDRS3OKVOn1mwVixbCvZ+kRnsGYsO9XxHTW7KJjXLsgFBU+1E4l
7dOkEMsRbSHwnexEj/s+nwNQdh8ilpK33EyLJgrgeks5F+YVKKo3qBud12FM+esy
atE0fbMAf3v043nFa8FLRxVq1jok1rDCT0bBNCQMt+TiEG9LFe6vWQoTPxTTKCK1
ccO0bO9QInrrlUbZvp0QAln4w1OkeBenX7bMHv90ivIfv5wkyIokLkX4IDVc5GyG
2nFlGU+lnLWLuGji8OQu3AvQ3AVa8Bp29kBRlDrtMQCQGRz/3sqD0feH+z5fJXHW
CvRrUnrC9bpN0aHjT9xd5MMplckBzDFAJDv+y8T2ilH7LUkxVu1cj5mfQfeQAugn
j88HH284x7SpNeFuj7DjZZ7n2E5R/na6gLVL10zGma0mIg1v9bt83hwUn14cBqsr
vpB3nepHYtd1wviwzQeE3DKoSgOpRC+Z9RM05SVKdsaIXmYPVVpYa8Y8wG430QBY
lmDDdeSQ6Y36argLyQXs7ygpQyFhQ4AAFgfBo7cZAWASqDl7gTEbZD1fz661fhP4
rkGwNGNj3XPYpL7sK4POygm+9akMSkjnRY8J8vb4I77/qYUL2YZP70stoZ8nYCYT
zx5ItmeUhZ5xrBugBFZITO4qIFY4JVizB6eZ0oOFFxX9aOR+PZCm+ajceyuv2zS7
bMlZwG161ShF1OwI7nmN28oH7Eie7UBXQCscdCAwrTV4sdURsTHShXE/3078WxJZ
ZE02EecL6NMpq6DVuC+KHi1NaVLy+yd+11V6Y9TGZyHLVDmdU9Y7QhF2Ash/LBFz
CIVRu62A6kaWR1PvKEdvSwTPsHC3XJB4ZyNQgajqEV3BAyn7uU16LFDoP3wAywFk
UdoWhpVSEhldPIgOa9T3Iyp0dCQ7im+T5K+qUtXtBjlIl0YEJ+lBOvaecl3MaUuV
yulwAAQvkZpi0f3vd/FGECx8zAYK3Ts+DpOPk+sHvwQ9tju9kyX9r3lrgtxFT7pW
MlkgtKExNqihOPzb3jPCAtVyLZ7hVI8vT7ckzqLNytcZYd0dKXClEX1NAqmeVfwN
uww7YZ2AIyGAYBGeIKBa3ofP7iN2Y1ONIaklvFPiclD+/nkZjk23ZUJ7UriVkjJ4
5Nt7pi9+nAxmJvQ03NiFLEP3iAD+N3bHmkXWrmcuUM0HvPpT4UmmJpDfEdOIEXEC
ZCk5GL/iJm/t6AnRIMxve1PMRs1Lc6XAo+T466gcV9eorsm6Ant1tEezchAAyG/F
w0VUf+pXYeeV3CtQoJRxC1KV5we9mxTgZdxy54tJ6gRzfMf/qYmpV4abOUrs3jrU
/fOgeFDkD7X8TkB9tSNNEgZjaPYEUc7/BITIjTCuevYGM7SluhLT8lq62iT+Vhrq
TEQv735wBqjpbKsh5C1rSyW09tYEOSZK+xzEArEDyoPqNgiarU8+pCuBMRGoMTPb
tf1VKgU4Hqz8SQkzLCDzZKB1ekXPaUQqxrhTLjVPzM3kI2nn4f+RDiS2YkFN/Ee9
g9Uj9qQ8Nc4NM7OAwTrSgbq6afgwJKnYFUFiPDDRr2adMKIRchOuEjOL3H3shcrf
3x0bsK4q43CGHM0ryy9KzQStXV8dv+rdOCTNPA3d0/M03yE6s++4d2j7jdsQGmbW
tm+QZ+BqdTfEe1JkR9Sa1EbdypQI2M4nLBx9t2J1KbjeIb8MxN9oFoxBXUMuMSHE
JC7Lfrfe6MyPRgTtY6UXumhDJOWZKMdeRJgukUxQmI0RluwRdAQLn836ECT4rx8k
SblTBTSCXrnbUDj1S9SeIEsb3xPTzRFoFC8sLwf/NGCw2R5Gcf9UK5Gx/IRG+4c3
j/CAbII8rMe4MdD0md18VsKLd8zN3j32rsslqe/uEOGqjxiwQ3LjPQ05XimFAVKB
efBzuJnct7y7Z4epSPNC+Yx+Un3uuIPKqazDJHG2EtnwiZv43oTxfknUNVtBRSLH
VPDOFrbi0nM6Aim6q+1Au0PGFhX5c1liCuPkvLA86uB8u7y0aRhujyvNdWiqLRVv
tziY/67uc8LYteiqvayEt9lyQ9VXtZNZpyxADuaUSrBF668TXo/Pk/1AfJMdMbBG
3y/V0RRIcULyeKUjOKqsXd7pjMBNfM7jJEcoXObxXe1ahFPILldAH1+T80gPF3/b
XcsDUB0rL9IrVPLQdeg3Kl7j0lee3ya0P/ur8tKWVIO9F8Ggz4nrWkYUlPf6W0Iq
0heCZ5ynNxYoOwwlS0Afn6D+kf4eeL4Ld6UnGeJXg3o0Fw7RmZEgmap3ZWqITBfy
u3+QXsNABfkJZW2M18rsJbAhSugDJ0SRiQBKHC/uldlhQYgHasH1Zu2JwApfzJY0
XzmSIVtfMNo4Hw8EhH9qzQdKxTWV0SrGmjAbL/8enO+PjbcZKgNFE9KxQt0HBUBf
gtrYgSmXGIprr989AiCLU4IHheGfTLdWDdlY5rtHVKIzkt9kF1sqDzhFxqPgUk7b
tyoLSDkFlLcRwSouiqE1RsuTehC/YaZhm7DgZvI7FSH2eCh3QOyx5ShcN9fGeikx
pm69uGWZgSPQjkFNavl+l5qDJAVIal6qOgWkTPHjgbpvUnG4tWdbYv9+Bs5p+4wP
GVoD39Ej6ya4/B0fj4Vo7Mz6L4oicfezciwHU1BZD/diyAfHEz1SLb38+tCuEGBi
1tRdIarLez0zrz3+OIUygsYnxTrVZEnhQ/C57Rv+GD4aybvdMTZ46R1FYKUURaSX
9GDr/Rl/85bI1Y9/KPitSWRClgykS/42oFGDRlPi3v3pEuGoVkiMWLXqrZ3M1Npw
LXL/UTxynqW2jj3x+rAhUA+6Py1YeIcZethVOzygH2JIwEBpHjwmR2IClxbGvlAi
AmfM+nel1g2uzRAOeo1z2I4m+1i+YF+RNqcZphCcYDkqt+vEXUF2GPkGMAAz1y9I
38LyhEJfRh7kw3Le9H3hFqvssHm+ZWkmWSpAaMku8pV37MusQrlETPFTuP+YQejA
w2kYeCyxe5CCIQnErt79Lylm1TPfLsrN79nMQ5R42zazjS75oS21S9XWAXlCv1Kb
ZJXsOI9lm7znun8ZrCIIbhhIqgMay2F68SaOkimEx10oH1/aNzOFd8JQP8g5VcCo
P52evLScHQF8bdBJxuD8e84jnpTgrHx7DIWY0cEz95U/T6EyPYM4f5HemJSxFxAG
mq+JY+1H2HLa7PqbH1tqPwxtC1MgMSPVxBSlefKFiaqkDvbcVx2ZP7ks9EEI8QBV
K0le1AwMTe0tw/I/HDD3K9Q3U+ETPdEkukDpLsqj2mSYxmIILmsaKZhKRyaYoDoj
DwU7hggUIe76x9PDraxVNEv97+EagwPh+47DdqYB3FlW5OOzYMhvCPEBO/OSeRCT
EsxOFZniHbT8Avm7barlcoCfrJmQBhg+0QG57GRsjaWtN83W7Q0kbK1nDQLS4P33
GeMR/Zc7mhVz1G/HYYAUVfiwWRe4jweL9K1LmtXJeceJovSzAb4dqBj31hKKHUg0
19ZBrqW4DawN2tDX7KLlehmQGl22h8TDHaedgYaAzPwavdDte3zLhp1Y6YDzSY9H
T31ygPwm468PWXyFHNJjedoN+3RSjqskCiE2leI7D5P5q/ohD4Kgf+FQun2bMpRL
cn5dJjQttiQ8+dsyPnKob2jDPWr6YYWq5bOgBgpBJK2jGrPL3mjEEg2qSnhXHNKG
bHZ4c53EKC9jDqSCsOSR38I1v5r54Vz46x0yuJo0APXCQqzvJN7rfj5ZaVHoTz5g
SjM9MIMKC5iODFK5zuu2WzGhghB4KQD9jtuSxe2OPtzQWGEAhqltRm7M7ROE30Iq
rGlo+LZNYyU0K0+DKyu3IOQYLwsDQavBmkph+XlU0sLBjSPiokCZ6Y460Qse/SYb
aQngWJBR2LjXMmtBYa6VTCqEHDPn3cDTIHZxTebXpfktg56K376m1m9GxMDYobjI
AprXamTm5VXViEeHdxa8PlNu9yjhh0jvvjvOqaoE2KXLjNRL4XxAZWkSm29R/xbP
fBfIBpREk8y1iZaoCBTqx5D9UCuO9RPSxn2WDetQExP2vwsEdvZ+mJFS+hEwj06V
nHIPwEYa18XJHTV9i6rq3htR0uDFbNA8/VIKWE2EebeTVdSLVGHhUlBbtHck5UUm
fpPmFpqfN3ED9UP/vX4mPbemPa6doXpGrZeqtlgfvkYECA/DUnAyJec8HNSJtoeq
mLuHKL8DgLfuXl3RinBxHPHdS7+ZCSUNm+kAefY2cZTDRrwd6GoRs5VS4yzD7w1x
1FnTLWA1L8+JdDkDPDC8GUzZQ5L494KVsmdjE8ZTxCwZKUwoKeE/+2aGcogCvgVe
imSXBj7DpdYOYWxqWzPtEEcH/c/maRQZKU3z4K7DpTHB4V4EHbsl58b3KYq4QvOe
ejUG2XGOPpZxpWX9WBDVTnRcSsnNCjGjb61VdqwOKSzsrfBY0a8P3JccwEbPzxcv
GeEt0kD9xHfnrT5GrC1y1VjOmbs7rizSQV3bKTJyidYywj7BAGMYx1O4LrCa5p8H
YBxPZlhFJdMjeXySlS3uij+8ipgCpDXImSj/TFMctKclamLURpd7M9FECDRYhbSm
6Z/n6qDYy8V2OSlDRi9hjIWgnINF7iwirQO+EqC3oBxpbpD+WpqbXzaMXfK73A6k
h5rQRP4Pi1TAVL/Tt0czQRTubexw9iH836sj8uwyITGkx7DvdsSqx1u+z1ZsUaeY
FIJHdw3EI0TVm7WMtc2qCVewmwwmUUTCkY9TtJ38d37RDdHJgc8JaG8ZmcU/r52D
tC9Gc3NAyWHRaJmJjJvHPNe5FOF0LFX9+rrztZ+xfID8lSB2H6M8LHUpp2xxRhTg
2KWO9ZjWUNgYU+++BcCY6uHTu6k5/nbGgjfziO/1E6fuEAacbqynQNEA/EC9kc0d
Yk1dnl6SgAfMdWG8tRYJTC0cFwQ0+ilVRfR4Q8c6nW40J9lxwNT25UgvkEm3mcYf
CLcfDfgP11lJC+huZYKxyhOKuwMWv2vpmB24CmOQT9ENnFK0siA0Zbo7fuoYIXvL
R59OjOibNc5rOQRWXHTBBhmGrrkg4ztLZH267YABcmioJuaX7Ywql0lpPrxGxT3R
mYzktEu5DWZXyeEjcDIAIfkcGqZrPG8v/i1SHlOl/LktISnzN1YR+rol+ajWC7Fq
gWs/NPDqjNqB8c0fFoeog0qE8BELhbNi40efCXWD15Oxrr4OWrT/VWG7jKIdMjju
x1mCqtpfd792FpqP61D+NmSZCti2+CJu9GUz3LIBDh+QWMCZQxXP85e+txmwxPCj
2HhxhEmv7iTlAwApN945lOd9y00GEIeDsYYoobTUma0ypqeaDEFt2MMxI6fk22jb
x4fDAa9OnjLuWg8U9A950CFTsY5IccCwUiJEV/61BpwY09p6OcFSeux2BB7pTHlO
7O3LvtzcRRao+VMy/5i++4RV95P3pWm+8ECElKcwVfHcu6do4IQPsdceG0fe4Mk+
u37XZjwHfXs0S4PLW5UzlK8h5LYZ1S42Ux2AN/veLRlNH9ae0k+iHKklKb5V2Cjv
aByJuhQ2QyKfUwkr6CRyI6knQxmamjpTDBafyozziNK2CD3G3Fto4IPiShC6OrDL
uViQFODYxiP1CygVyNDMOPOHDymBAn6qfxF2PqzJ6qywj5EZi3ZgzppEQR0fE54W
byV+LKVEHSUU9JaAp4IuYBNa5Wmj0rU5jpWs2mMbcWmXSaYC3ntVdoofJoAEEEOU
XypGafzTtQVkURIVmeYX5w0h0cIkZfy5VITIJl7lcIhGA1B+5MnPcSp3I1aZv1/h
gd6UQ4umY4C+QPg4w01ENCLIM6OqmjLsMX0fekghqEmJcBYkPr6vlf4gzzVtn6w2
Q1wJyFWT1X+N3GZvwUfyDZsdnTzH1MhTjK8iEQ8I1UHRh5zcB+SZ7KXzaKgmDIm/
gDbJdTbnEdMRmWMp1Nzj543qw/QlFEX0gS4i0UBfiFvv+KwKDIVJh6EqvYhXdZwn
dArYqc79wQrLAf+Nb7sS+mzucSUvK2SW+JQrXsV0VVoVVih1E+u6MPK5JXyD5RrV
zSeR88L/D/mrB3S1UwSwtp57lLAB12TOuiD6vn+s9LG0y8uLm2j/5xZA5yO/Xl5z
ghkkfiIunk2y/lwbLNWl54GqmB50VxYY3ey1xBBcztiv9Qbdt9xlx+QOuXgdibqs
Znjd7/LDQfuFx6jLUHZllQcS9o+dWJzsGqulWHx6wmUdpy8iqOIGyrzcK6kpQONk
qQm4YEDgExcHgGtA48VOBoffDkJGL0/GLQE5l6k7IlAzEizyF0wW4/Rc4Xs30Exi
WDggcRE54DstQCiGww2hb0EKnb2t9xhbfqfiYps+Zb60PosO18nOeX2e2+pEFIgU
qnWUtrmfQeYPDXP9MMc8C1LYdBJcNLNxEXLS+n4huLmKlo8QNJFre+UCnqygeMAZ
Oug73Sp30wwbYT910VM/CTVDnDaLpDIQ2V+H7pRtKPhRHx2r2A9dWJJA4M+W1rUP
ISmWLihVa2+JX33YQz7SLr3T+Q4PRB49for9BzaX+cmfA3k4dUG4cMF2+6ewuhQz
jatM7y9xbB/kDVK4NNEMSbD3Xm52kYTgtErbgXWvKIsrYWRKPY0OU6jX/HdCQuZX
yKhIVNG8KFeQhocPrXA8CNI4sRBzA/F2i0P6Z7aFayiZGSL/x03L54cWIRFrG6db
RqihN2lCP8C5R6ILRS4y5E8QgkrC8uXseIAovVS0CgvZkgXNZde86m0WRVGk7UYf
Z0TSYHLP+biITzfVrKAM+8twRhQRGa3VvYlUsDPnmOhkaYfjFRRPgm0xPlDIAcLJ
q0Adbqy3bZCfX4NhcXUX7xBaY6Pq3MVUDyKbodk6ksN1qfYJs64YCPVFswsGLXTA
7h9uPkH4exnxFY40aogjw/ZvCoYLTFALoVzciD+jHoyMkvU53S4KvChSO0623vi/
yGWpz6nj1l5mqkqgR2B5wRHU+8HyAPFuEC3rVmSRSmfPqbr3K0ELLJhpdJnJvXTE
+ccRY3yaWC6EEg57IWBj6es+Z5CVY7t2/UVth9NC9pnvrB317ygNVZV8Z/UbXi85
C5Ft/m/JGnOJS7r0gfMPp1qhsijhziMKnGTH6M/niXQ3MeNbNiHe43uGkE7Uenhf
4asnkuFVrYXEOZo+eL5b9GYMKjoHDhhFCq4OdMam3lNqaFWaIKx2U5zMswNeY0M+
a6xX7/7XmAs6ka8WF1/Tr9vV8FEN4qPRBkKMCEU1lpMMWOQXkRysZ29YYhVMHaUK
IMToXHxUckU8bEglRnb4H5Y0bEVGxc3W/u40B5ICcA4ujHxHaih6YYc72JGOXO0I
eJdTkYiU8xn7mg16bIKRuW1TU6g+WAOFDaWtHJj3wQDaLGk3KLvHlrvhZ5utvWNA
B/KFaOYfTaRAucGWoxdD/N3iYAQ2qlH+iePWNeEZyT9gvcIuQYnTiEP/kQGVLH3h
VbRFvwxDR4TVaFNd5dI2hPwyORjqu3OV+FRTfSRr+DLWfgrjTNG+S045l/TfXMVj
SvBWP2gQ2yM1QbDN+LDWtZ/BmUKRSfyZHhV3/Uf0XfU4auEQX0Z/KBn+wjkqWzpH
wBGEQZ+qgbMdM+/z6tZt91dOe5d4FZXMbjhSJCUn5bK8o+wrv0OakVL4xeYI/IEO
albZfgk8ZCPGhpQbEgjJmSqMB0wanhmpC/m7xgxlDklZSzdz/nLCXYV8lw8B0iZk
1+JfuVYvEYq4ZGJ/pnDQ9zwmMbWjd4Dwc34Ytm7+ka1BncXwHjHOL4zPMvjf/AMN
an3hEmuXsMM1jOx3aq4R4pPv0U2g1/TB3Va8T5dHEsnMU5CZnUc3P4ELJ/OtS48a
HdMExs9PKOtrImWmQ/swKeVFmdv35m2eCodX+RTCm+DpS0RAjbOndUwcMsofjJ4I
WinMgiSD8tgoZ/elb1WHa007obHN+miSwnGrPxegbfuYfr5x16KADislKxfXuthf
4LMF/54sCjoc4K0IYNdMMjAwtRAVw1zxQynjDrhxXrqr/TbU3On1y0UpxqYipoX4
33rGGILlVGldpuZLbqUQ2ZtuVlJh3ItnnaukCdiMHtutXHRcFNZbLuCOakRwiwiU
M2KErmIUOoD0fqSIGVOF9BcwYfIrtmkbHOGrgSHzIGZ7eCOibLAhsuDR2ef48JZy
sjm69NmR0hSZJKSPGp8ysdDr1Z0bMETyBeVSYqbQw9mV20Mi9l7c8v+nptJ/PAWP
sPQmfGTufyL105uoZs9jlL+6rKyDLAh4ZYhsApNcRUxH2IzAMD09I3sGUG0LVz9e
FF4rD6A/6G8lwi4/ISdcEJuZu2MZuK1TuXuX9rH5VIbvkDX01WFz5lnu8CxJqODx
6RH44O+7UBLN/WZIY5Y+K/nLFe5esA8c3qmyPihJ5EFKXJ/YuA0oPwXGDHXgobZZ
ul5r/uoeqql6vLjexnttoDi9uofQhNMblJx2Qhkmo0SGYFR5jQZ4pvST/Uu132EW
g01BTOdTDGDW9ayeh+H7vYLCk1Ao8WjEzgh/xaaXgzUwHNfpuxrCFSmOuNHddE12
bzwmO6F2veh8DrXG+o5ntBB2p0NOAUhENiHvwJDuYVQNZnOXOnM2yfflYhOE6fX2
S2LsT9r6Sej1mo23P50+Dm1iIS6UmRA/Y2ny6VAr1oTKowy8BV7x1B7umTwD9kZm
pnxEeKMS08pXcmtOH5yq17h6Lijv1UXw5/Uvtltr4IqF9UXwh3VrQE43wp7OcY7e
9NeZTinXGWBtPwYlfjGTlyFfIw5WUYdF4zOpNR38m5P3qnA5MWR+beN+57oI/CfI
YFVfEdKXVhOzKAUwc1KVPpKV24KyKHHFjSdXyvPGB/WPjwPRJa5qyI8jFBbgSCRO
5Lrn3TzLRwqYiszso6T2LI+4/vbfEhY5upQDkAoAcfHOoaNdwGBcthDwD9yvGqMU
TVF6AW+L74G70n+sCRcabDQNELI+0WjTkqqjkIyCUbRyLQZ7JGGkixfE4tfiVulD
e3p+/M50m8l56wuHurlnaxQh3E34BjtZ1l5d/MApWg4tzeW8TpmQjLk+qA9Nu29s
0ei1EaWTp+y/qQtna/dOOY2tWLc0ojN/3GvWi6z+T9Chb+1dOwbrHxWjWzDitoSb
X++dDIv7N5XnEfZTp2XRtWiD+Ptpjcj0ohy1bu5cPlhG+plYNQ/dMrvAVWFcTfi9
V8ugpS8p01HDlXFtmdjm5CunjkAJbl2TlWMOkAYnkxsVUNZkB2D0snMCbFeto8bq
Pm2OKCTMKpcDgJkLHfdI3CLh0NkiOAGxy0tUPbGK03D24NH4YKznXqYqPmtfJPs5
MO1WyIdvJrnRtLHgggO7617oP0yUcFpUL3+A6mUhZjtdVR7uBvufhCCAep1mKhbS
oIwOn9BwqodgRaqN9fUdq+Q6VJ6onvLvwdbIdCPvXqW/SjVoRC/kcu+TAJoFZHCN
BTVARYOXzv/fTyH3jO5ijB6IneSKyw275pSqjl6thdU+JNV8kj9LBTtEn4ruBtRB
P0DzFJ4FjoQI4o9xZAbhbj6LIP4F0tcP8bYFA64M5A86nCbSnOW/6XhqHdVomT//
wqD8PpDps2ZRVg3BDqa9IdQzq0YKSzcVbSdM3mPUG5YLCLXlInywh5r+3siaKN4K
TuZpOMPTlEFnONbp/8hEJ9VaP3B3y5FRy8z65XAskGUbxzVwtvnllp32ej1E0Uup
1vIHCAU4VLZm37geFB+7Dp2WpgtOZ/oR1cuOxO3siDRRzGmEet/FI5cZbSMk6nqH
AFSO9lsiC/GiMPdBIJyJtSGxcatDR4VwHx6Neq9JrLXOsV9whlyplsKRfEKoEHiW
s4suc5TS8RsqgkIpLBpyTbOs42X6M3RBITEj45oMLI8Ve0swxQ1/bJgEsuFSvr/x
tOsvyNAmmGBeJ51Y63ki2Mk2hy6f5ZPOo5V48kuA6j+ApcIB1Ygx4Ey9H42Flc94
UVS080tIpkcHWnZHp2GJW7mGqtfOImByURzoiU0zPqqm6pXT88PQOM8q7x3R+4lW
PG0fPFzrFmuTp4eEtqJTQxhNzf8SSKf5YIGa1TcMG2/E/7L1gePOiYwqyyzcpk0o
8Nr/Jqyj1Q5LleFJy/EYQPBhxy+By6+xiye+h21v8Bd2Fd8E+qmwFIb9J/5sbUwK
lny0TT3WGdmBpIpDBFuwmdWXmbpSyDx6cSG2dsrU0N7gMf2I4Ajx/d1ZMNVStdLE
qHA3caad/YYYPEhFTxBqD8CscT8SoSf/HbbI+f1HGJuJhN7ybJ11wkrtUTIq0DlU
zgF5tLuz93Dig8EEjh0UjkVdvdSac0YeMMyFImhXjnhLjDlNgTjbc0Za+0y4d1s8
94uLKTqFKW6cQN5chLrpeXCKccasNWaSfzXoe3PSrllpnGJnwH2OaELdEIA+mM9H
njrpTGrxv48FPggEHYh3i633a+CIsrwDAFziuqNUYEjQM6N9kN9DPVNNAHJN+U4U
TE1y83l5XKE6x6w4sDGBS5GbMZYoK6gJd6p42tUUuZ5lHN7Mio1IQekwO/dT/b41
/AyKXP3Ln9BUUMH46bqA0c05us78Uwsiuyi47eSMIr+/RbOQujE82MDaC6b2bS9R
vvecm8DWVMQWNIYrM8PQlr9+KiTdLUB91DIxiEj2rZxhHVvUvNWtGvCBU28jRsrF
tNTMecf90naEOkK+rHHq41TwYpD4A7kFFhh3OcFrgQNKsUrMWq/MX1wcRtIWD8sr
Zxg5YxQ9o/JHUVDOPv8ZGHOnfSW/GOe46pgKhZ8t2gQwysTOEFvQIejqBC2NlrPT
G3trCCGDJ/moY3SmG1jqkSTG7dAfxpuMiQB1iva8AxV0F00Vyz3OwlTucq/Lg5v3
1VZlPkabfEzhEaNY8pfe8+OVSv7Pl0lELJ0uOwPHN4yCdi9H2PDhxICMatQAw8Wl
sign/T1XEmDkHOq2fG2hcjliSlw3coAnRYCyrZDtbWtdl2gbUq9+uOzHDhdPpD3X
B0bt/K1Qta6bq8lNsrxLkqQmTQzvWprpKTxYghVg/avBCTb5Ohda9qzD2f5HGQyr
MsDwE4QPn4lvyX3LWYzUfeuPNUzgxOXps/Y4jOnSj/gokDJ/Mnw7+f+U2eSMq8QC
j+lUxWRG2/yvLCwL7JpHFzglJE2OanuxbRuigIjmSPVK7SuZ/JS6YXPfsQ6rWsKj
WrZKkDJqrGcF3gyL/ce4qTZt4OQTI7ezi/5HXz+8Aep1A0Cld3JAIz82BVTScxvL
u+ICc0JyP+gDts2jNAF9oyPEW/CVScKk9bVT8zZM01aszlI05v3t7yVuZtN5tJFM
0ScMMd6IkYRURc5ULaxHPThaLXF+oM8M8v2gnms4Yy3BNyeuZ81shwXnQzjfly1H
dX0qvTgqNexJcY6hWcGNuhEKD0cFAQfz1WtR1A8ypa6s+W/iGHofyY0TddZ1d8Ld
m9BfgJewyvxc8wF+iccqX3ZuQ1B++grguvv7ywvZ7TUp8kl8YGmAbbCwf90R92ya
7upodQjKvqz5h/BNjHWG5eYMLSFZL5EHJ3cByZkL2Gj7iFsXHjZS+Y87wH0rmQou
+1JfuC03VmKN2PwoZ2fBoLkD20+kBsC8KFf9QN4avOXVZS7UrRTFf3Gr6jZVa34l
VjdKP04lMBqEUcxobIpmiEJX2Gwr8ts0Jt6fgKy3dIV1Lnt1H7Hk9Hkp8yrp3bE4
HZzRfAzHbBVlJ4bWA/GJWq2m8uthFuVMA+FvHhmgn4KNXjDxjjcr7iwa47oor3rl
vqv5d226sci24U2Os/c/Fwg7VumKRZL04CsmzFClubhpWmH1FQ1U4XGNYfWbr/so
kHIjkl52IX2zDHxT+NIBAKLJ7DcNHE2PZPSEKqam4DlCp4Zo3cfeuVzjdDGJka9E
MtMT81X+JOF14xlAg5j4fLUp6kJWxtQts/5LfYB2dzw/KvRmUqy//y3ZFu/RvEhw
u0PdRZIDts7oz9T96ola5diRyst6R7Bit3SD9ZJlVNk1uNo/w1poXfep0zR7pBiW
g3HFFZMhZwaGhmlEopYmwHL0xbqNIEBIe+afi6oulgmm6xqtPvKO35qrMmDMseGe
yCJzFck3pUzHEfKIPAbyQGBZoqNhRA0alT6aAUfvYnqVd9THyALzMUu673cptIRf
g8TaK7bA8pMZXBNdX1cMr5kGba75vI4ol1yWkBbmMragH0h1ESJq7dAxYPnYyEZL
JTvhA28JUxCmlvt9f5FQyHQkB7gU5jRmL7zdleR1z0C2+Lkq3ypeMvoDUGZHzu6P
tSD2gmvSvPmOSdm2QW06XSBddPFU/jQ9ECGyuVUDGAtCEGvSSdMCm2EBZ04JDBOU
Fv/bjYW2eMBxtPL4D4P7IEeEAHBFXFjFce3OJEeklv97XAAjdZfOR8X14INM+E3j
lvFB0YYqBdjWs2uihZN9GSPBQyOKNQsb/Fka6YW1Q81iW6x+OeoAthBk1bTsvTQe
3yoVmtlgqox3NeiHcrl/zIwqNQ8HRWng7jkjNiXFtiALqgp6sv8oAJO/AxQzXGZV
Dvw86nnqkw8FLmvDkW/7lhGiPfqbmAXwKpjSb1asjTdIg2N/LVc08G+6jd95nhpQ
anNz1OOJu58T+FryeWLigj8QRO+xIYwvzhhepbmdrcy6HUDbSliN7L1IyPl3ix47
SXqHnjpqhiO2Ow911etQUtFORAASYuKNjCt5BMwsw5vrPZqA1yIBoujd1Fl5C0tK
Sr8MrB1ddNgmpHvJIXvet4vsmCrOA8O/PkxTcWsUbYfnvTqnmbXufbopYWkGdfst
VcRVmUwyZdHVWHkJIZEbZcVJE2O5nGD04Rt422I68rh5CdjvN2LJb5aaqUrDrkQ/
kj4nJNCRNfNNBaAFMIXlZrxNfzo3a84FNTVcqJojroEw5n4JpPdpmHMy6uLulFSJ
TwdwYlUiWUIhJFIQ4Z4+CXYkmGk1rrRmgGdL6reRVw5eg6ysXGEKXN0kz+nLXx4j
FOolGsc0cYboCWHnicm4LC9pLqXzVPXCsq6yNPDaJByMuoh9D/S2ir/dFMvRB4OT
Onac96YkedudicyysO1NZP8Dn/8ZBnb6T8/fJKFbWa/UltvsNUuGH05yDih1Q051
G91UzyWfRkk3CtgugJeYX4W1KMIR9nNZGPL7dwR41YJK4FdOEVWgyyjZOkgkCrpB
eQpqjrCla4Vz8jcauyJDuGQ/AZKqgAEmi0ebVHHok8CMSysJF2NLrICF5AzM3ruZ
4BbKps3m7nlMfCkk0WULNdiU1Njb4Q/A2mDRwUs+w/hRNB3H42cymbHECafS47AC
PgluAWTCDV6l2nXSnS6SqlGjw4SOdssAGaBQslO6gWB3EvsjkBiIZ/Eir6cG41XH
0I1f5bBrBmUhfKInlOCmvyZ6hFsHZMeUcC9QvyBaZ59v9SqhlLxZOSzqmg3BsyPa
9uAg3y52cFp+JHPPtvoQQc2YqfYKQgRiwm+z/baijTYi3QY+ueSNcifY5Aj4/vB6
RXBqPTimQ9XpZwuOeP4R1WB+5kDpxYpU/cFqu0gNWNzlcD0+iFoNZXehtSA2H03E
1oN3Ifd/8ZClJsugkyW7bEnKuvvOA64n10H0i9Ya2WNgTWq8wVosGMH82OvO5GbB
H72r0CIxg+Jbd+UuFG8UVxcNTfeuGBnts2fJg4wxtLK0OIqWqhjFZX82bm5+Y6us
Yw4FnXbVysQDbT/IBF1/t/OU8ck+v8MRvh9aCpSyDg3VCHzezkV5iFJyqbi+2AKv
2/2uHQfIts7dtbxpUrWQrfhy1CV4nNj3cy3Sh56PJSGNpM1yeet96ZAqwSYtw8rz
jC9O5t6cze2ter07N0CtxOoLPKyDWZaowfm2wiFpBG/ExFC++KDlDujaVZyrbuZR
cSpDZ5ftC+5TmNS1ic2IQt1ZXEo83cANQ8BUr7ZlEbLa5X4uDFjzJJyv8YhlHX5B
v/aAPGbUk/cz8okUzj2lzELHIKlMVA3/IzXoL7IbkQJF1aByyAv5XPMwvG5jEwZI
4gnKgPdfErIQ7T1lofwFdAg/voJnPMbsnep7OMjXFFHZyRf/BFqulCj0qyIIf0pX
YN55iYbFfZeZekh+v65f4JEv8sha2LBfdGluXRFiG6JA59S94dzKqTdQdhVXmlgO
DCmlp0mbIjE8zJFQVZ4CmsbgCHySgit7IeUtQ3eZ/betq72DrI11u591SoNOSmzZ
ZSnTGUj+mzu7+KDOxWgChPNXhdnNUTQ5FrhnAty36dK6C6CqCOgSvYh50SdFXDfh
RpyZQTnqaAyQnSSWfVxx3BHEXoBBrCz+KNmy9YS5yrFOgOL9J8McpQOfbdmlnMFR
kKw0T6muL8AB4zbFZipAD7xdnWWsXHnmfAEgN070nkjUm3xFEYpAga7NtMC+O9rY
llMITmFKBafDUNHAvMgEGJqU0XPsSTxpN4ra17dm/LsxuMg6N2H9H0Zh9WXr4f76
gGzqgLrGZ6KZ2xUnoxoqvrtXeLunWPaZP7BYM/AeBp4qvn3ciemmYUxddnqkBh6I
5xJbqBxVXA1ZUrFIffaVk1JrxiAoq6CouwxPq9oI3yi6v5lUFNTpMG/oycAxyyCu
Tgs5/Zy+vBRk6bJjmUrJPis+FCjezRmPkxjIcaQG9LydNXH2WuDfMQZ4PmH00pJr
Lwl947o8tiRR1bs55EExCZNf7gMXsD7UH/KZnzOMIggFfqELivsDNs5BQ0/bjcad
bWzGe3LCyDl3VxC4ChIz0NFQ4YKzQx0YYIc7+BhcIynBkIkHnv2CYCCFdONOjS/C
YGl7cXuYPwscnVvCRNkLQIWp2gDLV3JyvoewHUcPq2znhBf26bRYCJeFSyz/K121
VJ4g4Nc9f8QK7UoW5y6R0BA4q7LX+JlsYs6u6vNDxe+I/wzQ43j17UL4ibfkUHWv
+fdZ3GVg1gDC/rPkfvRkoQxIVxYfG5K0qSa4eSaniAz00Pj23YCN+R3Uzmv/cnXO
pnF6NAtbeciL4CKIVsjm50ZSqA0NfVlB/f85t2llnxE9R53xxCnoBMjGoIlTiyNm
UbTEh5/uEyIaL9Ggt11uf6FI46w2d9LIeQQkHnJcXc00aoLQIG6o3PLd4iyzYJLb
DRvAiD2b279p3fMdeEkyzxw7Mtzhzj4PhKkFUeuGCuxXcaQ8+ndgZbkKAQu/88z5
5XfHdFLPsFiyysEXToFz9tr4vbCMkHuRAjHx5I+8mTIaDLFf4Y/AISbRMiH9u8W7
qhZw2lnIlrED1TWLYyZ90Sag9zPm/XlvMIvUtyxQMs5HRMY2O+NowTbirK2kNxKM
cgsokixUbwoLpftJyx921sWeNQdHCJLkFwvbtAgD0SqLZ8DbIYNk0jUZUDcql4Zp
41LpWUu9q/mfhi/dk+kW4UlIL0XDgCwPTD9YVOFbsPfDC3FkcgnUfwuvtumYXBj2
LeSF+SleRSQIDMwsnwrkdmACilrk9jwu1k92JQise9qg6c7HLsyE4xAhkPFEQ/5R
MKlVAJtguI1KEQ+Pf9fCaQmbHY9nIJAmOSL3TsjTiQwk1ONcLXSMaV0cPxqdAQEI
+6RnCwPopXmsof8KMUStXlwltCzYkOq/LrSbEyL5F+uBZIetdx8X0ZtMcG7vrvrN
VSQSt7uA7uQHq4vMh9gzoUkEcdI7Fs6OsAjTtk94yAsZ5wFrxQii9MdMLDvCeShl
lw+D+VTo1SKqVdmq7b+aqtpH7LwXQW0+OXfY+sMyUML07IRHTfqAG7tB20M9ATx2
qVy2LGCoeX01MJA6Ipw6iAq4dHToCUvwNB2FJgZGrlkD2PO/5zKTMZP1tU41evlT
4V+pRVYYuyAbbjWYI2tY5zdNkkKDpNqYp2uREHKi1l8QKwI5Ffagi35Ier/gYenY
KAaofp3BaaWIgHgKLT7z4fXdcvPEKUzCxspBE67OKrnlmGzhr+iMS0jfZSGpizme
DONytslW4ttMkbv+Vzu/f51uvaGrRek5edMGb5MG4qIOUnXopNkX2albanXaAimJ
+gVQbVpNf/oY+f9vVPJJhIvwgaawvm2ey5yKVi3dT66pNSZBRpE3ktKlR2K6/c1v
iYjTbeQ6OWOwQm+aslN6bAHYTnGJUifah1M4VHhR7VMZR3JY2wzebsgdp7kKEHGC
x/VJtsh5cLPd5+v46WY+G7jpHM49/MIbFXed3F7zmfD2YaggpwpgLIfjQOmYyjhJ
4z4NNZ0soENRvVWuevgrc8njXtIa/qWlctZNTKNh9enF+/uKPO1tw3sKZ235Lids
jzPzI90MR20Cxz+2QZu4Wlb0OtU4IfgCmN25HIHdEI6gme3JugwI2+dUgVvTDDXM
Wo7TDy/wab3JdQ2dNf9QgmsBb5NRg2lXUfC930YDH91qZ2iZ9gyWfZRemly+9PKJ
sPuDkl39Gd74CY7NJuSjQnkwZTlJ1Bep7Z2fMVMVs9ef+gtC5Q7nT13zn1ZIjhN/
iG8lsJ4ZrzbM3JqIgiVOtNgNZBKZJaT1E4HBWdpiErkTD7U2uzvKh89W9oTNb1Xg
bUkBoBOhUrcrnPlh+9NBK91wko6p/6iVTM7Bsr2L1XO3gQUOPPjpf1EUZQvLtVYk
XMtFfsXBtPETA9CEssB7ArLOkzcf6hKdsuVf6PaAa983AIS/LMZup7yP2oz34Vww
Z9kUYpc1QSAIxiUAduWL937WZVwAr6DauYmmsYJ/GlNyqQUhljukZrmnMpLSVjwa
Po24i1WmTJhpFRbnc+Km7TRMdlv2x1+OAD30g6vB254vRBbhrJ7/oO5zYjLrBTQF
UgnIbDR/ZXboNNUISbwn/VJQiOUOgMaIX0bKMlrfU4xg1meHR1uyj5pm3RN0EoJy
Ya7iGdqugq4KRBZ3GGMrXP+pj+827FEkwBa4TD1GkTe47edbz5E0ULo92JvotLBN
fChoVVLcvUGksyAO+58az06WzC1km2FamYTDXmna8XqINsWSBt/KVYpUVwgoZMRC
IUt2zJ+KRFn/QR0vMKXVx8QZIzLdGSYo0cEiWAE545XMKHZdKHSv2qh09IF+TjIF
Y5Y5LHiUBmAf5I+jp/p5bRVi9SjV64+dNFYYmUYnzPKNpTOLLs9DdyFC9nu4jLeb
JZ0MbCvYtbxp2OxUyXX43qGtRAOvvdFMaraOX1ADGcqbwBB8HUEdITN90ZJPEcT7
vgV+MiEvxE6ca8ovg2ynBXabs4KCVMWlNvCyYu09duOidbFqqqNIroPoc9Zi0oGP
/UGykQJIZQ8CpsB7Wy7PaJVNPN6wTTELltOSkyv4ATZiM0Ym9S8To9artfmBMtZh
vXLLhE5NNWidjVd4G9KrPfAruOX83PwY31yccO+xIjrrmE2FCac8lQWQLQkU9+x8
OH3+qy0SN3WiILWguik6z7sJl/oYNGN0EDQfuulRLm6SYGUJjGUNpNEPwFHNr9FN
0Bw3QRw2Iqnm7HaTwvnJ9ycXlTZoxAedLKuCLIDxoefbMwBluWPP6xja9BIFEdGq
OVsnrTk30z7KDWeFrcns1wD8kS96kB00hILSo7QZCYCoThw0LPvlZiFo2DZc1IU2
mc/jzq85B2IU+ugVUtRcN1FVf5Sf5FljmiCUJLGLkdDuePOp0AznaVm2T6IIHB6F
IOCKB6rjMADuvLoy6iylBxumGSQ/cA5YhJnRbcfopXOXyBpFUTzik1q/Y4JyMQDN
AkqymduO8PqMdTa8hZOC2ru+Ffb9Qd2tn+QEf+0aK5UknA1lgDu6MDaRbX6dQ9Q4
X7hAaglvLfqXXhMOv59FHR6ISetTscfVkk27aIs/wtl7GuCUi3Q5BCLF+lSYJ8yu
BgxpWvgwFvo1wOiKO2OckVG8P8HnQ1DzWhuTOlSGBE35Y4yBc0vnSUUB1ZGbTSbF
XtV3Fd+o1CDYVjJkT+TrkrbBLDC3eIaahLuv61xYyzqUf0AyG7THpHGmCHOdnhsl
s1v/sc2JndiAdj5/vZzbkBciKjvaMxOD7LPgwVCYC9Rj6hjdJeRB/dqBbMxp0T0C
SQAIZt8pEYwbbOrRJcA71SjSF6uYIHAT3EQySKaQJz+hPJqjhNb4pRfdA1modUrH
gVkiUpzh7JC5W3nAmhTxTrOrG1SHkAEZwQEMPoWAOUtatgyQYJKXZLOoCtKLq4+2
WwTSCqUgvquTNEgpBvlhm5AMKFeLkiAwCm6mUbGOUo+//PbBwoDHBxmdIUq3xEnj
vUp/vL51RoVvgMcMA9QSPoEDYn0pO8qcqCBGeEl98bqDEIqV8Q7JRXQAJs0XvQC3
gygbUlNlhJrYf1eeWfjWTyQwRVQ4g2FRRzQuso6r6eHPOeLypQt+q5xAfnaQSRV8
6RkqvP0rhufIorW1RDbdOfdSFQfC5NhzoyWMoCzvKAfrPYbpIh6iD689HgsCdVlH
aSqmrgtE8tkoWiu1ykReeWI7jKz/jdLuyezAF2r59DLdKAk+8Tac9hdToBcTJ78a
2KUelmv8ZNCiSkBo0LlaT0JrYOU0o7WBP2BVrmQsh6GQ9AxAfBZJwPS/0IZwTKbe
SjgBEA/a6sxz5LsAeW3YmK7tA0v0JrWS/dQonIYiOEMd5DWC2qeHHo7NZX+SC2sI
hgxpXVYgJZjwJgRNT+XudjRnsaE5rGys4hdv9WwjJ4BqhSZU94nhljwmq6ZlPLgi
wPBkqwFeEkQ33z8TFn8xWxSepipakBNWm4Ow6eSTL8DgmJVl7Z+8AxSdYzt9sje5
/0GJ0RFwwSz+thqo+9SICctaU3ivjLf2Cs2BFcPh+/mttOP1JIypKCqp094qph8k
CpwslYwMeacIhvKtBfYlxQwpXEACJWXLQLURx6i0yccVj9/tkoMknDw3MczRwgJX
hQgI2qabu3G+tTuzlSq/IVcpbBhYN5oFI4rzkPeGK6iNIkAWue0IMTbaLTsI3qtK
VHcZDngvccTurvbe9sOsoagtr0pxUzkRCVGwxGHO3/Qi6o9wssgWnk+x/TgAlasZ
Dz1HhfYOupR8ZL7ImcjSvpkfWeK0vzdYnjE982rf8YpSYievC90KmSB0ysgbAt2w
KPcyOQNlgVSQ042pEPacqjp0mYOnR+fuBM8f3aFPP4W53GR2gj2Uk51tHGVrwOSS
SpbgIJVasSp4IA1BxzJMht9VgiEtPU3G9DB0GFa2wu8EcnBr2JDsu2F0tGy8vprt
Vkp5pnONrKpcTImxtaU+/WtK2By/ejb1jSGfCnlJ2P/C2vMwtmccaCTW5yBLe+5Y
f60wAgdSrG68NaXg8Xld+DM0jCaWR0EqrDn+Afy23OajYqEZ3PkP1CQa/eiWy/T0
eW0GAH3LDbXTL6vl5pMWXWXfiY4ZOYaWJHnlw+wjs5Wwxqo8FxoCaaNFmz8XzJfH
iojSS/rQVb5hsBZchPNT/apAZIcVekBbxxjSyOLh6tRncOeI5X0IC9EJGmkbnLd8
Fyg46/7wK4GLj3OEak4dKfsZd4cGBm99VmIoyH43dosjiK/6fZq4Blh2CP09OHuW
beRmwtulIkCAuozg2klm6D2o58ej+rz81ZUWSIlA01IxXfhyKPuA7fLYTxFYebPX
xx5SwXtnyOCG2oW5p1TDPHxbwMAnSAx6BasHRZZwLZYLguk2oNQyEAJFKql+F8zC
cMXQx7RNQlGQQovXDsLk7s5C+60LFXYM9mLhql3T12bcdVNeUpsrTDzXvoGQUvti
CiHkag4x/zG5iKkMeKY564IH51PQdwCpaVqltFlMO5bFVj2R7DCjTVXf/omp73dA
JqOIS7j/2EkOKQ4SGUKVf4a5wF/fgzAm0jvTFbD5a961Y8kZvGu/hKkQg0C4Owdt
trdK7zfJlExDzAIaDwBXEw4Gzkv77nL1m3UUMiiECQwuAjQaKaFRvL5SbFhBCIi/
jOEMnrDYWyFj/jJ5G5BT7BCxex8Gu7vwy7w70NW5BXxMWIR7XiNvNWgxpjtmDf5+
0tn7JTOtI6vbMlhrp4adyDnvv+tTmH8INbGuKKv9OeX2ln8arhfrms2eYLgVN2uW
QhlxLQsjW6k2KKJcZEhmFDAO6AGEGf+LaDYugO+OcuCql6Fm/QTiUU6MCGNrCUm6
JKlVmS0QK2afOKr0IYForvhoxgY4x0TjyyF5l9i9AYFbUdw7QT+B3a8+dRJ/19Bh
bjtDWbV8rGeb1WJH2bd5DfL6Mn8q4tPGAdiob+j/G60hEH1VSM0rHDIwLr2cdkfc
CUDU4TRUzvEqkeyGakqb0psxr7sgiaNqNUNYsLC5Gz3lOjnTBJHzzFwkSOx8OwZe
TtJqlbrKUvWeP0btkE7O64e53glXnhTji3snvVv8sj5HLZ/MjHhMT6+F66bVH8zO
NFOEVA+abgxcWd0cNen16JcT+nmRD8uXYzQPgvQcdB6s5UoTdsigBB2p2TuyMmgi
j+twhYz7Hy7w5L+/hGr/WQeGH2LEPa1o6LISOobqCyuKXNguWDrkHZ6E8FEZbuqP
+4liW64Rc9ISmHGhWOmv+b71FazlU5momIlaq3Ltr1YuoAK/rTbm5zHLTAvcMLKN
JCiW4nkNF0RyIS6tR67CutkG6aUW8Sc3zKFwzEYo1kZvLd8mVvxOC5pt6t8KacTp
iIjU4qQQe3VrHFhAZoUf9fay8Z74UyO3e1FtTIr4j+dbnx0vM+fIIsKvpryu8spn
zdkZ23HxCthysncrKIPzjNn+4eyyQoAL9il/X9ZFCDXjHwwyF1Wq0otdfepIXjyK
SrEf8OK7r6KlQqAQdwg0EFpS4L/J9u5wzCeOrCRQ4Ti78jyi2dwgV3kN4W8f2Ek6
lFyY1848EaXbpvlocCBBDsI9eq4C/MpE2e8dnmdkIEEr04xVZdLZnI5Rdx6Ngyuu
0o8nHV1ROikXIWof4oTgWIR/h2TBpr5tgpqwZ9lFEMFR2f1F5BsHaHIvcFBX/yDu
qRmCm5RErlGKc6nfxmLvnJFbglAFg5iCJt36u77A0aJlIi/gPnm0zHSZnwe+aVPQ
CjkpKc3OfsZ78GM15wby7HapynkNCEtj2SGeiPbJeMf3YEY0BNflxN5iY7CQw9FJ
cLV9kndDoo9/pp+EmsWgIexYDPMQErVzLxodbl8rfrtvEVNdY7iIlWWSDageNRwG
NoRABWg/b/Vn85/sJ1wXrNFiH+TGui119LYlErgWaDWBHK10ZLtDlMmiAH7CGsHm
DczfkfbKmAJ9u35GmT7UofdXQ0cRc1AOAAxpEtzxthNfrv02zOx+MWHQuxQFbtq7
W5MhKn4XASTcmFX5xhW4x8YSd6dCGhPUFHoQNq30xFIw6XN/XvrGvWLsTl3sCHrg
vUa4vl/ZqYjIiRSv2AXWqVka1mj+kpQJgQv6MDiuGjc7wL+k94DmCjiA9dsumZa/
WKmQ2inCYDa+GuIEAMRgKLZttxm47CgjxVuKgd4CHISNJP7e+5yTaT29Eg5ZKtO+
y0yh7+DitZkuR2/PqPtSjkyNln4e6GLhuQu98Gik46e2k8g2ynqY0F4KEqECh9vO
ZDipPz4xFZ1ypT+Y9Cy/O4PDVn+6A5+H+lNp+8Apd3JX0ZCtegLWEPTqQuaOvwso
Ve8vS8wQ9othEFZERqy1cZ01Z+RA/2psd9jn97GTLIRWbfy9bfeFrhB4EraBWdE6
7BdLZl0/xsYC5XdjBzRSyrlsBVkf4HeHXmMsrutxUfcEPOV7JfsGMLWMSkB5D884
v2V4qOPzcWynWrvPRwYnsTc3GAqG8OFXZDZpbEZxvD14hyN2khQb4+5XMh41VJHG
p/xJo0upmuWqNQmAlm6wTBngh3YNyzj2pVn+YEgcxfLU8duwggCqtM4nKmT3XtDo
3HVYUuvtmat061ZsSk0mpaYsv4s9vRiShHXWPFXuhOnkdVxeC+H7jDgrfXVJ8+aO
i+m40el2h3WVw7RDZx4xj8Ggzm9ppVdqgqUuk94YnYsrTJNbdXBp0v8dIpK7iVSr
GkNSff1pP4hJtpFSA97tlHPUYVqLgdvlkuZgQqNxylsfpHV8w83/3EVuX6nksSH+
++nB7HgAsBgwVDDxkao4zSqhdLMHiqz0MBb3zQQ6SysidUv/4yVAe2F5ebCQo9Yi
vgDDN5CwdXbU6b32dyGEOssnTm+4jMzaNrVURVe7r/YGX3Cip0a+v+aOkz1FQ1As
EQEg0kC2pwvsSLNFd/hfLhhUiqjt9XagBSUSyO0UJ7TiBnwitYgtFfRjbFw0srrY
O8xHBQt04S7bEMXxeAdbWPLMGQE9sRp6hencT/9XD3CRRrnqW9Sb84K00X01sq7v
pTFUEwLpuNNvL5gNO6Dwmg/EZE1+7KnMKNc0EzpKwWhr9C4n5LgffvV/G9OyKuvU
BBzmb7ol+0WZQitGzFztEOhuh+zWD5s9nJrDM73iJh5V2TfXBlrivOzAMCXyJqKp
eCzxv1J0raDrbEbhzLYiIgOcZy2EbIlrbLr+9jYgNX7UHe1IlFdf7oalLESEScZ/
Y5zuVRNXLLyyT9jigGAcimYFcv28jWoQls+pZ3AbOWALQ+OANktudJdTwkqo1Ul9
lnFBiLUAC08K2oh009qCJBnljYP89hJs283z0a8x0fHm7dcRNWWR81z8oVHMtLMI
BKSUxVtLTdbtlpR65tnELGyfrmfXu5V4OcKvDyaRtm2j4zC4tmihgLuADD41QTNi
HxuaGIXAlzjk+RSE6H2PBanmh12gx/wUiZYERKyHxC7gDwXwJ3hyu3otK/bemD3a
40pbSkHshLATP1qLQr+W+a8C27KeZnFIbquD+OyYoVjkbEbAIBC775im+S8uLWAg
7Bccv13kdZqiRYfmKSMhZML2+r6yYXn83QGudP5QjriBWV87uVucmtmawBo8WqT9
himyUQe2qjL8uWtHL1TtlhJUvz7FdV7XashoesqGoKqbX7VzlC9AO7yiz0s6UrgS
aZYWhmsVeH8BeRvZj+tbmFm6lSSb68De3DVEHpRHBMw30OC4x2N3OCZ8sbJeDdru
2Gn12jDkCz/DWU3jKTWXuqWil9CzW5AJfXxQjZRT/BsyoXg5GS+U70UDU/7h1Qzf
x6pdQP0VwjIqSXmh+JYgBKoozI//OvsX/NczuZRnOM6CD6FpTdnboke9U00gF+UP
rKhsKyPd1/PoIHinTEAQAv/AQC2wYN+aJSvwyT+kvuhaaxBgR+1cWYyrTMlBETLO
YtcgUyaR6oaer0KFlIKp/g+Y2s+39oSdk4hwVvLUr49EBxHTy4TTb42D2X1LaRK+
xhM47DvyzD14Epkaab81WHA+DNgDEKvRWCWE6x+rje2Hi+QKjwDO6Ri2Mewk8qqs
p8JyMU3u/shPhr+bTAdpYzfDCrvk8I6+wc6uBLte/z/hTKf14zPhxWkjKDTkLVwO
W7HHpqy+BRA41qgAB6ecnNIYaXiq8u+IMJxyxpp89s0l8bcZI/F2RhsxY2a7bscM
gI4pTEIQwZGftZWLACELhxfAYl3f1S6PM1cDwIOnTLQuf6V3r5eSOJlwjGYzQKIY
bAUw+3vTKP8rWEOCDdf06sO/xZq/x7jGwWTdG5gmVXSK6CkJ38aC3e46nllx8FtJ
WF6cgW03G03D2c9bEmDZd9qo3KIoz3ttuxcyZ9kn6y4KSrDfo4sBElc9/cdFjL9w
8Qn0X/ZqjRpFoRPZPhO5awEWDXFXc3ZvjyMRJXpKv7ZspfF9mN+Ceu4KIqfufYlA
Dz5Btx8lntYeGOD0XJEExoGpantTULvSByYQ0GYYIC3Ug40szVSbHIMcbJB10MxQ
smQb8uN/Gvzamk5FYpGrcHbWLZ2wINJp7kukn7rIA83vypWJ184l+YYLQw61TWwe
JL2QlGd7xi8d1fEMvQinr7l6NDQt5uqYdZ94B7D3+BSkoSBVcsu45RlhsCi8BPw6
JpF52YO4srM0/+qQqq76NR9mICYseyho2noy2hvv4dU9xiMKOfqIOma08aorJ6Tj
MzSgvd53aVx9QMkz/wnX2F9w5YtIwEmdQBvMB04mNq+v/IvrM2AgvPyjYOo0W2KN
546ymtsyApSGmfIUBdEbfs7nvRdqKvdSomhhfYLJXCXmds3XdYcUTQPHNoamU6bj
cAvx9OakwFbW8FKhRFsqHoY/8ym0UX5UFrK6TPdYR6MtlPj2YkH6SE4gLoksuzIE
UCsXZwNHYpU/DKU188VUanDj40jyqroyOTLyYUp/phWLDgIVtcUE424vXoXeGTVN
D8JicKpTzPnO/OLiD0zkjqBxuJXD6FdBG9hc+aaXfWYfYs+qqrtXS4zvAlqf/45B
Z2fn6JT83U+cZQeSPkLQRoO3wzN6v2leU8UT7Mnm1UjtbeEBvsNrCdcDBPVeitRM
r/dr5CP4eOq7RAsUFh3T3rTYv1FzT8P3eJhTCrp6OQ4PKekq0/qwsxWbUhFh1PKB
1orybhF4t/syV2qCJks/Hi4Z/upInV1gSJXK0GaVhRrl6ZyGCIa5Ewoc7IOPpHN9
ph4Id0gYCp9vd7l6fmp3R1WrAJhKNB43bPBU2ITszi2X2igiB6VeB6h8/WkJx6g1
CpKipCh1EGIlxNSvRtFp8fOfiBOBwVseTMVgS5kn6C1JlU9CKRlnBoTQyDHxPLgO
TZczNPKw22ouFxAj+UTg1PyRluEBXqlGV4S4PUVFC1Li5Tdh98Xr0I0JXKpjHWb0
G7ixn5/DAxUQQ0XKQyUVYM6lD+zetgZFEgo9rSuUoFECrarZLkfzewrFmK/dHTKk
rntYVv4IM1ytleGyo484YM5AXzTrdruMnDwMZpS5IznvmKisR6EvsEmxuvl/9Nht
mRUjGHNZ3PChITLGPrXRDfVef5aBjz83LP01ShG0FAa+2BIO+biAIj+HO9ibedXh
w2q0bDKTgHVoENgKhwKP9tj7xA4R2veYpe/DqIjmDs6J06OH136fc6DqDF+9FxTw
Xrs55FhUc8PcSwQMJepSExOs2zb77/y3sHsK6jmPr8cZUDfOxKTSJOSXc1OOjUcN
knFC1mSExRubtDeO8H0lI4E2S4BjbMI3xyc5qGs+UcRxsa0gwb/uplDFg8cF/WQ3
u8mdtFsHd63ArYNNzM8Qu4rhH5TDWkNAhykhxTn/oxQGtxyoOStCRhXOKljf10np
UPREIQYmAwQvJjaoAzXFdUSvNpPQTVIVFRo1pYXuWZptQc3H2KTM0nKWw5v5mENG
Wd5F/QePOEm9P+8j63iGIcCQGVnkqvhg9R/eBrDjSedKPd8kKtf9/Y+TMX5SlyEw
gK3XiLHI6HEYXgQlJ71BZXobjGRkU758b+q+0atknawxY50cUcC4VwW1FDZ/HbdD
TLWwFzOLknRU0BhBEvDSuglEaWx1i5F4h6cnKWNcHP1bsxr7qTQNNp9b4+8lWyTs
AjfoOUiX8Crrqakby4SY8CYjS/tpwntjwMaiVXAef6fQU79rWw9J/w3W8JqXozR9
RVjabQPLg2sqHfbvZoAFBV4pL3hfXILUNa8QocquvhbUz4gRIvDAYfYV6JwS7/lB
3zwapefXIs3j3wQokG+YDarRmf1H+7C8MykaAOvTIm0s2Gv7sN0qibRtpvGRy0VZ
z8vLq69t8eYqdbsK1LIpqPWqK4m6i6pGA19tWcIXkQrAjcthWv5QEYmKta3npFre
SzUQikXbO/b4zmOZun2TEq3P+yV1UMO/dNi1R7NK/zB0sCCo8i+geKWNyj5qmv9h
0K1Yj+NoBV2wNYcSyTDNJA/SLb4F+g5dudttlpePjqRuItzVurSpuHLNWvGOoR5E
WFp/NmfrPFE43sHBqjQVJ2/eOFJzHpVVgDVa1UwRcROJK8G/U2S5iktrpvpbWbPH
9I32F0UNGR6hBHkQ0+TFoZmSHXTu/KgOpsm0XXOtW7WfEHQPUO15zf7XKBFO7Rlt
MHBrG8+seLQzvU1mGloWg16Y0fkTzoRl7SASV4Lun5wV0IwUoBjnfbkNCdk/fYSR
FOhLY/znGsrkiM8MkUP3iQn5XIsnsf1nnGro36XwT6745UBTRtNEWDX7lVJVhasm
ZkeQXMZ1tp7L1vBdejn+NcQ7veLUh+SdRgtDav4AYfXcHGYkNz8CG35p5mDvz8Vz
ZnCbU7teYPn9y2clRo79HpRraRW6hUw+BLQWM+YzrT6TEWTAH0w+a66+r/+r5et5
zvOHzghlMy5bCtvGs++8z+sXGi/hZL1Xy/h4oVyKCNLqVA7vz1BENZ6n4rp0hiR0
l/rKyG/M5NLlEBg2L5rNUh09DwjCPT33l0kIrkga0wGjzk2vsQOrHUNJaNjEQbvE
Q9ArvegpKDu1sTKbTqdUn5bYoZeL+y0PhaiFfxxxPwmAbvWLz8MxZWIpTExvcyLZ
DSCmi5uTvk/46aHB8MPWyY1dQtlYx8b5HZanVy2riFM1Xd+M5h9MQxvy58Guj8hS
km132JJomDmJ7OCuCZGjt2iz2TdTt9fKyzYlXSnL2tlYyH/DCtxjQZc525lfxwns
Ctk3ecMpeDNkyCE6x1gJVz0m8j9o5DQNoOvghX0crqnh8YWJdSIJ7aoG5Kue0dJw
R2Y3sJYbifdnhGFqoR/mcGxLlA1ujNXknEDOk/DzWRsH/WFkw8MI5tjEVlqsfqTG
1ZmEQOn5lEGZUm5+ekZgeLDBlc0BEK4R9T5b1vqeBpaEn5ohsR5/l548Py50kjzR
ZR5Q5I6d7DjGtA58c5gIdH3lTX6RpTb+b660COIITUlAZmiXbN4AHlrAdaISbDXq
bgnAg+84D/Z3asyodFBk+Pm1f7OTomCQFxyHKVCPqDipPwbh8OQgb93DbozyAdS3
lQad/M4+Ntc27Y3GDZAmmvQpTfLZ0O0zN4H5YTq/AMdQx3c/1q5o/vUVpi2rghOo
vZ6FqBOeIcYrH41xrQKO9Fn6AnK3zYb85dMC6PvgwAHprb/SPJeSH9Vox16GrMrK
KbHLbMwSFjU4lO/fVztiJErzQ7GYz1Ft0+LdDEdbgyC2M2E42e9zO5tfQs7NDvZn
GFvPYMfgv/n6WTjQfABA9elYW6W/E3fviP4j9TdBemSrZfK/r3Eg7AOh23DCHaa8
vw+fXTMLGwnAL9Bn5q5dS0dSvwmcv2QLN5BQkJHnSy/+V93ca5kPEpG+uRqUiPir
/dLuN91MHL1TkcplvahTE2e3TKodOF8sdd8A/bXd1+CU03uPmyKNajQCdYfY7t4d
N1qGGtN31oqXQASWWEtDvl0wYB3nBFLBsCecCE0/SgKWlpW7wqcC5SC+E2Vrk/OH
w6KUoiNpcAJ/iZdNX7PA9ipPWbVl+jj3FK+XkHdISLWVuYdaNhxQAVKxxbKO5ATz
VDgRZHCfiguiKCumnOjqiT2Y/URHixHJK1f+ucCXRq7szGVIc/eUMmRSOYF5e6GA
RU5zrYQspfh35Y6b9uCYpJ+dIHEqxg3gbGfThWCEnTKX+zjPFGuMwuG8a2gJ2bLe
u1YgKHoQJyDatqCZGzBIbQSCgMyt6SR3anjA9t1AFjVr9+S53ZMiFAPl1GQ0g11T
BWoaprW4Oz/NTjZPegJ8gGUFpBv9x68rtzSFzbSJA0nAlpLLu1EmGo0gXbbhI7ss
DAV+BFuOCbqj8AFJzaNuck7ruisfT7dsZhC6NZPLDTVPEZT/0ElJ4U4IKkmrCOMP
iuWiFg0LvxDsfCgvv6HsAcULxLHQZkjnutS1/22yWI2Oj5zEszTR3g7u0Si+WNrQ
9Z64Q/yRY2+21F0CguuCPrAXEYFPQ6rJulEMzDa2AcU8y73X6Rucmvo2hyyEtEEK
0mIozOe5Xa84xxhpsLVmFcg342PYjIxrWHPSZ+PRl8NXbCR4RBNEt4r+i/+chnch
h0BN2ylj/HFe9QpcJhmzcdFIZs9dNKmXmhirxyHG5fXu+/0ZoZVrjoL0d013ZlMh
gHFpy625OOULnIItepQSWOCp3S057T6YrVm3nJIaDUwhRG+02GlHRhNK8ihU2D6s
F3kF1QeQQM3PbLaeTzbd/JsSJ5pNSIOIaBGqPekPl9jUesVfWodHQSKss5mGzHkg
phHfdfRpPDT/NveHHBgSxw8/SHwXGYlg3AYdPG7x45Zbx8gW4neFdHvBSYoFYLjj
LZ0Mq2bc0UNLzJ2+hp/pg98I28w9LnIHmmeke1SNzrNQVk9j2viRXUeSv3cDFUE3
8j+JXFP5oVBVOp856/XJmS6WoVZGePDw82oybzOFm61jutlbjDWaGPrWk0XVT2sR
TZt9G+FelTFltTBnl9gDVPMs2qKrhCysDyQcGRtYeieTX/AOcDjUhNwhC5ei2V6T
ULDcHiYADesgpTNNUj8CGZFvUyMnZMFKAHZo7MiKF7Syv1crqgG8as6rA8XKt5l9
vprtJnXsLCzaGA6IFoUViSVJgF38tquFocmt4gskdrToQtIeZLoEKCeOroRPQiUq
aWjiJ5Fny4SS2AdO5FVg0+iNACsqfrEnVWi89ggfohO40g4i4EAXmSPRgfTzAJij
H4nnZLAV144IxvJVSjBUPByweBWtDvWgLSeSxrDnjT3amQ5iEq0wGKAPgUQSlqbM
2rxLS66YGIZ7hbogiAKUt0fBVdVlSaLgiZyJb12RjCXTAjqYpjHuvxcqqMCYMaDx
MXeu+HKwRiUXKqXFQfsZXq8TGiCaQFfX5wJkMpzVuLV8gf0HUeyDNaz/a9WNA8WP
TNyuxVaWhedlbCjJDI/40m4xg7WFv8sk7RDO8SWDMa0C1eFIISRR5zMjmmm8augH
pZK9s253t4sy5GezujkkBKfDouFJgx0gZXN82x6e4FC21ocsAJKMCc/vQjXGl5jh
j6tLG1MBEuAA0mvcHlDML7lXou0zgFvsMmXxfIQrzbm2ZeIupKfi9dwGuI7x/MOa
9bb9sEoECU9GJcaKbub0gbU5QURooidIojgtkB83jIFEiz6jbeIOx86cj6znH0rA
Ds/QVKVKCJnYlF7M2zH69NH0CF1dXo/aXKxqgMSb9MY1T5URGaILCC10+BZ86zm0
lYCmpS/mMoQIht15Z01kE+OUvb3eRzN8I9WlkQY+jAu4zJSCpdLjIDhtcSczjU36
AYWymN4mA1THUAt6CgQKly4utMFhA93WKB9Jbbv4P58fFfWkQxkxp0a1uFjETnxY
XyWZ9siWrScGBCMBdf4t+TMJI4gnsptSVmgQcM8h4aaELKH/0YOaS8CxILQ/Vvja
5sCKnAXBs8w7+g7rFmzGk2Vj4/R1MikHp1exKU6NoyhPhffYjkoECtQjjoIXrJub
VUAdKHh8RGkd9/+LTCdOEVFpu16zwPltWuw20f8OsJOGR6vdomv1IJEwpltwWZqo
ThaNWsW6cJfZOArcYGLIsI3lZSQz5n0TWQZg9IRvxwrvK1TUmASVzTzM2l691Tm8
/cAO56M2jNAuOaesdWinfhFZzGrut05SbHrYvUTPpaGnO1C9rftxj+sG5A1HP4DF
Pfa+jOAW9lQLlBJ3YCnpFDfVE0dr7ubYu6pDCFvq1UiqSVZa3ZxJfJT6cCyN7e9B
JQAr15ktGKh1VUBS8m2w/X0eWHHiKJjHAa40ZDb+omtsQXVH2v8aWeTPWUT2GXjZ
27xmtdsVzc6qqOD606a2vDslHIYpPMxaU10d0sx7woB03edKNYKLTdV/IcL0zSk4
POZ38pKEajy6KwIVNbsMH97NoNf3e1+ojqoQofzfDXObHO5lJ088yJRkADqG8MjR
+zWijHGPusdz+ty75dd0auP59t1oOk2lGIcTgvBhdVr5d1KFjgjGaj9S6qpo6CCZ
7W5+bNsenVrIhUidSQMDn0K9/FVh4j3iCfi1yn7ZhFlDaTswcjyBzoo0wPk3i1hl
i6wlhda4ATTQQOtDHUwq32pFvlowKl0Uhn98ssETWY5aGvid1ZRWUNg65W39ynJZ
jMUdetkU2nm3Vs8brjA8UKfdu6xcQajqv39GvWi+/tZWeAh/PoK/AD1vVKtTyJDn
s8BOriqsZlXkMcHOPYcVDpp5bj/mnpwN52mAJ4paH2+H/7bSiGlXNmk6kzMaqWPF
MqAz0/1HMJSdWaD+lyZpRh64XKM/ca3lWeVu2OvbAEycYDjIVY+bbV04iRHMN7dO
Y3LNwOFCWCjhbsQaK+XWSguhsP5LAF+ckpK3saMXcHoDYBfy61Jzl3SkiRsGJQgB
H0mzhVhV9oyS16J/Df6hh/EtXTXXoqCrDPYT+mdyg9vLAatpELHoQ6Px22Xp+XCJ
ns4ACnwUAZfPfMMF33qudYSuFrHudt5vg9m4BZE6yXe3IvUA0l1QZCBAsikrLKq/
mKSPpYCeUoLtvcseew/NuBl43vTmUxgyWYvjS3nkFz/RFZd7ujO3yBKMfdSY7nVW
v9u7U6km56Fj1yq2tdU39rZbWYJc8zRnUeQ7Jn2ncbcwVsxhYQqtsqJ9RyCcVqZH
7srydKqCckBKNnRQV2Q0fYcshMUX4BU5Yy9RFVu6VGG+szgsStD48V93cbCgqLW/
ZrgVvSlw8MWmguS6/1nqznGbre19gYLbNlzz1yRKjbG+MFTwmIyYrgi9uNyumNut
od/Ng/OvlLPebEMSDjtoy2h9V6P6Ow7DMo9uVsROrUj4rY8OHK0FB8MOrzeXn96s
kZThvKhfU8Sp0nCxvGc/SvoLJSwW1IJ+/qzBA2aRJ0dfU9y7Z4MPOhocFWxVNwOG
/QPd8n0yPDaFN3D/bG3G/NUr/fkRuBoJvkbs+BUjBLpnqoUgQhSaNHpTSmVB7Iy4
pCLh3bdVocDNfkZl57QUiapxqRLlrdFRp9LM4vxQzizhQTJyA1s9OdjEzOyM6th2
V3NThO5jK2OCBv6rkQAzRBJOONnvkuKDXjEpcD0GBtg/UAdR4eSfyWDjR8oPGIQ9
UtUYiG7RTNYFvzMXMK/pM3k//z+mHhDp0LqcIrSdAdJYpAFYhGoYBZrB1hZG/zyk
8YhxYcBkIFajrOSspYiGH+BimopZuF2oleTvDGPJkm7JZW0fBROBDnAua+1zLBqD
qH4RF1ln2SQmZC0n0z97bhcEyruoyxYfAzjuFzzbAbwBon/tNSr/8vXVpzeP3z0G
p6dqeoW9f0Z+HKAlsoZtHdZ/rNyxh4UvemISBnl/dZry3xeLywVVaim0EOanDTvN
M2KpuBDcDqi+OlK7Hu5qqVibGKIgHVkN4bgkXOOGHDKd9pr9FvuFKSh1AC4s6+wx
6TV6i00yjsAsyUCYNsZqjz/m0E0HgQaHNyi3YWFFz4nQCgy1LwDzY+11ICmHrWFz
8OI4XUoLTMLWm+wSmhHnO2npC5hj+tCDAtfSwzHMJSOG9uXmQTkaP5sqwtCzcQxN
eLY13/qVRThGf0ed4Ej8+U26Ctvxx0OJJxxAfwfdFGv4C07oKiuBcy40+52FxV/q
RZ1E7MRgxFnwtxhBjTD1uhEMW9HlR+dnxBfHVwHGLSXo6CM0xqQkt1MGBPRCD+qz
vT/kz+bRdRHneZlaEtJR/NHzmUWSvKEiyUrckg8sEdz8UnxOD9K3Kx2RsyoRw2Zj
fgZBHJjLGBbhUVtlfJLzhvGzlaURPG9w1t1A3vVSvG/GAScYpSuMgt875ew6dxM3
iyEHYAuqOgtTl02tc60yufMxUHOSEZgJ+fzqkNrV5gRG6HlGm8zeklHL2uzkeqzj
CCqgHqYaXL0dYMyEHKrVJ/oHXikKAfm7hDzjgzBMgeMzvZhKPN9SvMlnOXn7RReJ
dzrqQ5CS7J8R/teplPwUTvraYExzyL8upGLxmGYEKsPTT6CdAhNtW1vCQDcMXkTn
fgjX22iwMZfV1PgkuTzfm9N7endx6jZ7HRC7ww/zmi3VfML+geyNDPJdtu419yBy
4q2ggwGSHJDUE6s2QH6juo5hQeUo5zx4N81XpJ3ggd+cVaDrcjlCRXSlXcwlYGbu
oM+CY56NAOCbQU+l8uLQE8dzufNcE+S7g2OFTVsKxbdaqhEtwbyQ0zQHvC42FV4U
bORArcyiOdxV/dCTfFHGH4grEQa60/wbcgHCSYuoU/DwIDqbPsgYNAq0IX4m6VPH
SGOv6UyvIht9o/qWEbvoCLppGJDA/fYjX5hbjq3H551DvFM52k+8HBOr6BYgEa89
DiIxmP7O79oGSmSghLNVhhCqlQXPLzNyOaVJY4alHN0muHp3kqG+X+Z4XqN+u9yP
2Ubpsq/YdpA9jkJ++0hn2JFHhTf37ONN1CQG/YIVQtdQaF0BQl7tnR5kn6uUH+Tj
ciX1mPnSJnfywLe/hlC9ONunJbFwQ/M05WirOhKCBpGurNKvyz+L7J/fOgjmqhtV
VduGm5b3QXRK9Y/pRcuDZSBDzOpfw0YbTbtoX0L8shKPgWffUcj5uSfAnUv4yvn5
etwF8tL6il7GdgUHXw/uYmenqCvTm1VprBA1x579JXZ2JuPoRWC/TxZiwFIDixbz
FrVZCuF+Samf1cJNJMCA7PoCCOTYRrjVrvSvolKAF141EYevcuohs/L8Xo1Tqpoq
Obh6Kt0DVOc/8gcZDSZgHVbjVKOumqA6LX9RlXX7m8tQ68CqWEe+wfWLv/yFYaGY
6ZvXfmI7ITXNUcYlnL3kWQLx1KwEnJNdi4N1FmqvOALfs0c/dpSqCckGA7KuRZNN
K8OwV5b7WI2F9IQUo/6NUcBBoXsAjGvSb3moFk1EYfrDFD5Khos9L/gv5pfuHgbj
3T4SRqyRN2NtMdtU5Rnh4CB5rX/+EvWYZ3Ag4mwU6vN6HL3ZHdEhJe6gNKyTQfAz
/p0gJ5ZgX84boWpqbMqow5OJOj/V1VrqhloJWA3wcTPHe44YUv6PJ5oW6AqtPki6
bfWCZrHXTTGSP4fwnAHnfnhzq3Jh//9XSPQR0y813zuUHuzZGMw8GmZN34wXoxl2
EwZukzui1YxQx7eSUlhGw/9TpTDs/NIxJbVZLwFYWm6PtMFHRWsW0bXx17GAvXH4
3Tp1v8g5ZlwywMDWo4QeYsRol4rW9ttPdTsRdd2CDrDGpbjNyKjVvsrSvJWi+lsQ
7BiFhfVe8nGRLa83c7MIEo9Vm7N38i5ed0HkYQ1lDa5H5r7H4SkQE6s8e2rJt1J/
ztND+qFsT7Zi1ZF3LYRtw3g2Ouqd7VCC6/GwWMeoA1090xQ98auLwzKqK4Gx6Vgo
ZSeUZChbUfGe19LGH0L4E3cmYg4r9/2PfPInUbQTTQEu23wdkddk0WDhbZQkNzeR
Ole/Qc2Wjy+gFacbYSA+5xa5t4dfpR8r3BMOVRfNFfp/x8s7d6glzWMKE4y370j4
mksLlHXaYYgwyyMZPBDc3a+Wm5vHW/xM+LrlXivcA2RLn+8eRp0qfczozapiXodC
RzUsw0/aGQyt/BHbKgBuFWp7h+iNcbyuzgh5vnpUzco9fHil9vl2ovFcfLIxrRPt
i19cqsWVA5lclYp/fWGcPeasafMfy58b61llQwgvKhSc9fDkXKhAy48+db5ec2H6
lXPFBBj6yJcPxXnUFFf9eExlXnKAa3koldgP83NcgXvhfZNamNMc299eLhCoRYpM
KcnxCLjyl1M/dVXd0T4MQ5fXPfXJQ1dSpzOmScjQ+RZ+TA8MjQh2BTDEpR3qSHtt
txtpmt6yqY/tTvGMF9eIJeKcmSLeEA1YoIE/iKWb6xvLz/1vLuYxCzEAsyMEB1rL
avUaRK80bY9td7RqGPh9cU6PVSUWqDnoORvTqR/Eujcus/0Hw5EvlayZ708w564T
ae0flZ+zr7wCy+ejp6Y/3homRdVPaSotBcY8zYQviXekhFCvgJEXg7bCS82Es098
MVAIG8sqLrz/1Lsj+6RgnBrY/tq0Vp6sCkuggHm9eQ8a2zmGQaqU/rMABokq1ZFZ
V+BjF52pb8ooOR3Hd+E6+mCt7uJaTIj6kOCdZBSPNlOJ8LPngOH96OgnGJLaTiqy
t4g2wCmqGWmaGfLZnQdRwdNUWhUEm8V3T8ObvYX/bsZ4uOa7/QkEeskNBNPzn0Nh
rfiw8Cww4WpQ2or9J5lhyBpvm1W3morLULcNAl9mWEuE310oS1Sbp97luPq69TIV
0LTxmlEaa9Btt+ekjm0o3cBXht6AmbmeW8WkRSv/SCzaD+Cy2+q/LSp0rr1m10y4
c1urF9977GANd9vQ9RxtFNsFHqfT52jxFrsnilEkh7VpwxIMafUcr0HFqfW282ID
KbDUX6KcaAymgnOOMY6H6+6znCJnZ4bcrNrON+ZYxR2vrMLM75EWzVH759wrnRGp
z8dCvCoECNOn/lCZhBKh17O8Texdx0W0FBIrVposvmRIBK9GYOmItGHnQ388wdJV
jfCXa7oSnuT0W33QOEeambAwf8qETvfnpDjvT/RzQ8YlXYzWsKFSXADFzVbVY/cG
rTiDHpaCRpbX22UljdaWkKTYspxnrAv30I9PJe+UiR7yTP/mDs1BWzPL49dUJK7C
dfqEATGdRDsDAhZtFlrXkkpP+4yTwEL+lNpANgOyeIHhRIR9/tvnWq69xx/2Zxft
82DTn2Ak8Qq2txtBvJ/sO5B/KlHnvjbhbCLNJyi9Jy/oI673C2iGg5/NMSMY0UZL
B24YhOJiHv0ECS/aGGhYDfnaym1vUNv14bJ5L+yDr02JTpHol/lCl4ZZUa0pYHh4
hf57qxCtTryZXw7hVVnXhEj9KKRdYI1tIyfOskvLMVY3xpYjBR/v4HeWWusLm0Rt
IZp8bC3v2C4cIhWOBJwISvvWq4XjQxEGwDNTCh1uslBZzduLtBIygWFy+qPr9mbH
gtYqOmSDrV00rLTgzQeG9qLvWFJVjdmmNgF8voBGAyJ5nZar8seS9JfNBC69OyAu
+NJq6Iix1l5hOaZmydGXpCs0kzp5pLRD2vmsuI6QM9sq8AVlW5F63Td1flFKR9gL
eun4vuOnZYKOfPeIFx4dU41B+d8fDvkGmLkuujCagEKdo0o7DVCIxXawZVb7JBiL
kOVuDPuN4wmVxBiEMkKB4puWCz8d1p0myJav+5HWVoC7TGjfEbviBgZEf2cxMWNk
LTxCHIVZjc3j7hd4xmPSWR51CRELy/mkennoHQZjjZGaJQOkJ0PzUazoOJpTGl+r
6H+hE/wCOyjBZvXwdVogxX5Gjo+VvGF3kIlHInWoOWIdx988pfNx0y7pinQ2y3Qq
wKh55f6yczCPqvlRzHGlYKkVqzFdAtXbxBDZrcaHs5sxeq2NAM3sA6/tw8wKUU9E
fRLguFgMIvWfqDC6LyxJ3pxDrhnfvBrKuinWI0C7MP5eR/F6E+o7r3YNCpKQLHDr
6/U2ZypqF0Zf0wJ84c2Y7o3U8kSC5PlH/yvU0HF5HhLyOjjcssOX9HQyufXKIWjT
SaQv2dsKVSYs3mlgyj/OW9Pa+wHrmqnjgEz2jzNYazuu7Ze7XO8f1rZsONt+5Wi5
RHqD0W9giOijbpXJ5200Cvpy8sMQKyg3J9W/J6VQ+U9PEm4VE2ChJHrjrUgDrTAF
JlDGT+TsIDOxo9pcI11WXciODCqVWEl8svgz00Bvy0pfN2m13eOjEzGFE/Yk49Hs
jtG3FkSvUGNeFLWSgH8j9wYiofTfJK/yLKcAahS+h5FRhslZZSDoiVz1aNyWHsmX
IeAfG3tX5ZgoOp0mAWD/S1dP0FRdN6cmNR/4efaJQKb2EDq4lL+cFu5DkuVK/9B6
wGoTKeyI45l4xPtPgoQr2Ka1SBlcv6xHL0IgJTs0ejAqTVYlsILvgkeVZvHfEiNE
AWjg3Qe8CgHVilK6Y0k8SmjjvcPqjnhmK2P3NKKlx/TxNOAyyE9cFJf7BAdhvm7B
uTCqdRp/UGBBDkEHjha9zY1gh05/7xg2QcS6Zj9w24gWx/vFqY6zAmB+m94UJolV
wUPaTqqaBHRZ0UkHi+NYNkIbu5v2mQnvrFP1xbUbUR4kahDwKPXHshv5wyjAtAyB
LnShI1FwTYa3LF7nb2MGRpNG77KxMcYcIaF6UAIvTqkKWJQuFZy1t/zKZvlCPTxq
NihdZ2z7DnVLl0LHhkae8yKK6PFhw9cy01Ls+aVyTxZsIjyegJ2qDU0E8CYFTipV
vK4Kh0GjMRIqvwVICtJEb9rahq7ZFmIr5LAv7gEjvXFCHHfxRBI/hBqS2BESCbvO
GIrp1VAgRleP5LgDYSBnKjan7EMTPCRGSMkpt1EE8XE642N32Zp7QVHT+ycGWrwV
yzLeP+9ytlxDmZxeuUl1otC/dJdUQDdjaGHctd2ivQv5MpdDOCwN5/C3UGEa9QdC
VhZ4kte2mT3E/wRUh0Bac7msABXkhG+Oa6fDHAS87yVC5uSrdTMzHOimhRkwesDo
TC6mVpDnTuDHw9SLlqSpNR04KgRFVs3lw9nIvUBRkwRTEimVCv899Y0GYsoqTX0N
P8KxzDiSUOd2TCTeeOIBp8WroP009LGPR9adc9xiwVJRbnh86JSQaVXKH0Gc+sou
lMsJiegu3nBLeEfhMJPASmV/EGlK+vlb/+Zt0iyT/XAdyRWrxJd1BJht97Vgw1bC
CsIZM/H770X/ppGaVJ0wHgezu/4ve1z+QnKmGkILC98kTA4Gi0P08cyHdZCVunvp
KOjZ7gwdp+ZWiMYPM/UczaDhfdWaPyI+00lrDUtlZf3scnuiafVlFGd94cCRZ7Fl
KIQuOCSUZ9M1mKUIhjkx8bFrabVbxVPN4nZLaVsUUXNZISefM9juwv+4Vx+guvBN
5lLFgEzqRQQk8zJmxPG14oFiROweClxw5xDD5moVDE54jPEuWzKg76Y82N8vY/e5
6sZGGRPCTtHaBdodZsZJNycjfEkLwhfdHf4aiKii8kSkwYvhng+cpwM6sZN77wyf
DY4tKSWCVKPq2fcpi1VEUOOW4nffClHJDC5e11gil9za+nQ+mntuUZEJ3h7vss5J
AkIuN4gE1OkSGwwnAF53H5D+lZkRef/NgnFnuiGdKhoBN6yi7XmxWB2jRLXQkDKO
w/K7EKBWmHfma2PCkTqpUKZZCs3/ZH45cbjDVkXdIKX3qnrLQuzdt0SLP+FNUevh
XN3RoYz2ITzEyT8FENdJYGm0IgN2E1Jd2DWvxjAZV7r8C9FN/mlmimV1wo7pU0E3
AdGBTdORNBPAKoFt7e4paKPrzRR1lboMDzWt9ig+3pbltuV2NKM3cqQVgH2X6rmE
TMpcndIGLs8Q3csvKpIjRoFmFRCjgTSlf8DBnxmtc/VpIzx/sONsAmiqr7xIk0cE
bh49woGb+fMo1T2RrYPqIG6LlyDpVtvyGhCvVpKjFWeIx2yv93s1frGYQENhYt2S
1Av+A+FtfHoIZgjwx+MTvfSpGpYE25w7G/54HVzOK05L0Lk4NuIp4Ags+qxyIe+s
V10flgGsALmnd3gTQaCQXyOesiDBr9V3UN59pAeT2rC76kdWRGXSMmyPAIa2SOnG
xFrpX3P0B6fwlViXlqQfgaVpdbpgIO0ZKOeUT432hlwFjD4yxH3KVHKBc3KEAPOv
xW/K533xrm9yK1Qy6WEiVKZTm3Vi5kVYiAF+gYUxuTDm9wHpTL+qJchnDxXhQXDB
3QYN+3ME/yMZcBQG4MiADmTJxX3H5BBXvB/ugLmcAfp4w9N3He41YrcppN9EJ5/S
DuszQ2qbrCFjh9WudSt2NTlsUEdLCbVCtdkIBXZGMzbbGX5Eufy5wbqDQKg53IfC
NiMeADPAc+T9xKApM8EbgxANHhGZwCYY7b22HL6Rq9DviBptXu3uQ1hOcs4uXHsn
Zuuv0q+p/kovxTAOo84bcStct0a+f5FTXwfh8TCZBiV6FlhLXlZqVWb2HwxpkOH8
cc6TH20GC99OyB3eA/wPWzFP3mwo9kOvjFRWquCowjFeG6TI8NU0014eaXS01YP+
5D4WQumfCHqFdoKhg9cFp4VvlngKcXuGO3m9oN6ofYgBBFNTMJcKyCRHbEBEdWen
TlZbYOKIVUJpR7I6ZRNSD9JAEpN44Vuz6d2sJaL4AczVQslEL7zivpLVVWUxFrK6
LcXzaG1RonjTeJpnvP3hzcS1gsNqFgy+V/bO38Ckv/S9Syii0h9fRmUFiHGViH/N
NAbRnbgluHDMvumRzCpHCjCi73wnhYFbVe+oOLvJaa3ZZlqb4M3duzeRBlGzDEhT
hYmaa5wt3qKIDf4ddF2i4MWFyMr/atroLZIngUyC/AuV8rdKmlG7M5ZJtdzJW4u3
YLpR7UxoWAGvQPMMeztX0K3J00i+JwqoxqDi2aSG+HGAolAKQwzWn9DwT1MY/sUn
+23yFebrWOA/GL4q2PEbAMaWFzlBT2UXYkAaLSAgp9AexHBTW08O/eH/JJR7OYEf
UoBwuKgqTYYiP0gY2cJdUn+T71YXvJ0cWT9VyMUSZrEeii7ZJTeUA4+oNQl5R8VC
ZR1sHVpfrRzVP77ilYbfZaHRSwC7eRDFtInM9QXBIhGLW/BVeU7DHxKVlESA/U/m
uy6NDXXG2ZUYpXNDjmFZU2ufMqitt5VOQwg7N/Dz0XnbjZxO4gz7ODLZ2015ZAx6
cTvWx/FBYPtS2uOF92fmq9iDl2fOwyH28DHkR/sE4gucM5itZ1xe193bIQycj07t
Pp8TjXuFfihjLpyZNVhrQHnx9L+354DSBofnAbyORqK12nBvw103txu31HXuHY57
3XHPdCjEI1C/TgSuMQ7TBoLwqetcztzJ21gp6vR76MfqUERlpUuDzq5kR4iqfSfi
fER6SXQw41CfYEKvsUyP0GLQESGig17mp+oVlIxLwfhKmU4t1qAK5g4jHf1rLfFg
M9ayaolmhRvPBEm0lrZXPxn2R5rBhAOFPpVLVBThmmCmPMjrJO6tBSvkrdfyVUrN
wk5DEoIb0d7JjlC8honNFChwjUSCkd+Bj5dXHW24ljtYtOhGSKLm8wvCEnRDP21B
z5CD68jfR5M+JjNpQJmuzSyKcTcQEwzkE/OxXsZ8VwRPzU7UTjY62zr8Pecm+0Rh
q3pTEhxoqZG3v674OfS5s+9LGizdMLQWFE+cZlylqDMXlVXfThqure8/FFdZ4q4u
7bSbY/1faq6piYoKk/UhlPTo+vY4RhrC/Ft3ukajwMnlyyc0wF/OSiqfaIBCHB/Q
bAK67X94tal/iwame0K2wdCrwLZGNVi2T5ywzMGTDFiES5UjbjGvSR5RQLpGl8De
caEbNY4ieqMHY2w3Vk9+B+bR/vCFh3GWwBWqrHDfBhVECq371tcp8YH4DiioFXzd
5208LfqiyU7882p4pGCk5qmvk1ldHHaqhRz/CHkTw/6PUyTFJ81vyJtQSnkHRZpN
UKXXtUcRpk6axZWFVxmJLc3VOAsNcRFesNnpuDqW2L/V7kbHsZ60hx/6k7ujPlj6
uap+hV8bYAMUEhiQDcm3xb39ZEvOZIQc3+sfpk538t8EPL3jhmodQZhWzXB8JIyP
V3tKR+BlIjW6mHPLLcnEwXTF4YlD9iGzUsnXRhESSh7Q9I/JXpMLtTvJckshPxiE
+QzTt15s+6+oWKZrn+Jx6Ccvp6fI8YuUfRYIrvf/IuVBUOuGhpdhjuZzP8KcsejK
D88vwekKTeOq7XZObgY2PEjlUQtt38/HY85U5TY9piIomcAe2EZg7rQTxs5q5P//
WJYGYTsT5X0r5rW4NA9ya+wpyRuhQcSL+LwEC3C5hZTG/aWTyPJtUVhD14M+Jat8
kwJ42BCihjSqfL1PLiPnhrpcpyUe8w+7LSUhB5sIAu+JOTkeNpNouq6ft2KWi7WQ
IKNwrGM3aaS0w/PxPg9ZAUJ6AG2vXlRf4mUGMjItVFaOWYeGTdMSkPWXaAqWmYBZ
TdwIFBtouQdGW5OSPSIWp890xVAIdjEIoTkTZ+tRZLWU4sBPSX4t2tam//iFzkUw
1QpQ6GC6rxqDv5Zjr4t0QQeScXdw21vOTTjGZZ/t0VQ4NPAPaMWsSCXOHB2Erj7T
e40vZGpyCg0fkR2QzBOZ9EcIHW19vNEukB5OvZxkduKJH/ymQgL3BiISJ3dfDu+x
gDEd2ps4dFs0iQdUWtt5rtzEiHr7bqvYH6FqaLHV20RNYAsju1WWfY/45eXw7zSc
IKDpFget8oGrOcZqHnVciJ72Q/kJqwOfYkk0+83UYihpL6u0dEB9Y5w4G62rl/Ua
ukGbdhUDfsilX5Cp6gla5Ydfhk1NNcRirQOqFKxd7rG5ZO+1FFGb4yWKAwYA2/aA
KzM3jhAghUWgwysfrMRAd5HXlEBcCBcUc0WwBkWIG7ok4Ce1VX1Lsga6i9Xto8XS
4WyAfcKw5CcjXiC+ej8coResBe1DipjIXyFajeIZPCkkQZd8pZL7UY+ll3Ky8KSo
pNjoRBOjz2KiYMuzYB06ecQ9BM10pblOJjW7aECFeQvScZ+pmv396sXrhaDsoEi5
zxBsU/UddZXMmSKsVvjhXXNxwp7blnnkDGCDygALsmUHG7g+RPwQ1av244Jg1s+L
DRaz+S2ouDAkXH8B+l2KRETYErATP61S7ssQIFNOxENMiTY4cPVJBBqGN4vNWfuR
f1NAEEV/1IfyyCIoRkJkV79pqw26QSjyWglvA92QzHRbI/4skhlEzsqufMXzf1m9
SjFhsc4YdAnNTxL6bzmT+xwpXNL/iPyhj1xVs6C6VqbIjBYWj10grNe4Ji5iBQan
IPqyiTzFDOgUg1i7P2RH6GKSqHCWaL1k43GZJt1F/A4D6p5JL15H/v1iOCqYtrgs
RiYoNjSPpx8PyTuvuKDjP3Dh+c4vR4njB2IdmNcSVl6Q5YJoleCCjIr08AH/P42g
Drlx7tyjSpbVWLpcGDweJ50kVB4p2zQ6fD3B2CPFhyK6RsGznuWcBhFZ7jRRdjDT
u/nZsLW+sOf6GtBIu18duDmcNz7f7p9vNYXzKqt8UzYpL613jYObD0riyOOIHNCZ
F8SgUOsjYk+99ZJXugeCgsbIsEK+orMj1b1kgUt1UB0cpXcFSN3pKKNdP8j4aW4u
sicJ/GrDZjJvgZqrYPvMx8EYiZFxW5ncc2OUb/NOdHh9iYy20yWGioMa1OSwHktG
vZ6O7jf9WMc0wF/z5pISmVhXpWijFEuOIP3FgR9oLn5XcNTqE251D1osI7yH7xVm
adE2w9xPj+PtyYV/5e1wfAxEfDODYTSVUTN7HY1SAHy8MhdnGJHBu+I8clM+EwdF
GR6NlI3JkGZ8BgoAZ8dEEDAdVbBzzNaOQ3qdT+OymoFzCMWE4Wm9wTcWh2YSdR1E
Wuw3sARvPYc3tPLOzmoAh0zJauyL5hx03K+t0c3CttUXNscvdlTrEJioTcDIB1v8
vhiM3qEtaYpM5KqzQmtChw1v9vyuW8nyIbpX9YuCaiS8nIAJzR6elZ9bYlZnaAKL
SA/GDHA20wSCwBmWg/rH+XhRUnba408v+7eyvLH/+Aib/wMqmEwsfg8hZgrdTJN1
IfajJDpMuofV0mc5yA6FpAzvyB8LLqxUJr4ZPPA/D0NpitYf2/J+ja9ksIcwLg/p
Xtv4zZY+NcRXImAuAGTrviOtH4NOpgmnBLex+zSvWBOb+UO3CbxeUI9nor9TOR5O
miioj1U1BkTM/sPv7xwFZjHcYTpxqxspFYaoGsExpJ9hGXP5+9vNRsauCv14DZK5
+cF/Ks5/gHdfRijC9KfQSvyZEWv4imd/mV1rnOUCyP78Vyrij2D3yxrLbdnNtva9
KHFeR8aRHn2Ow3qOJz/MfCNyoxZ1qDEl45KlR9Kh42u5MM0bmY2aLetx9wSWYuiM
X0kDNLl++auM6OASabZ+Ha7JB7SZjgIso/CY0SMAo3u5ykHvCMSGGgvpMxv+avdg
d9XCuk7mdz5sa4ORp8INBGgi7b1xj0o4ACAy7YdIlsXw7FTalo4l562bADZZQs9O
yqyqDsmV7ZQy9W4MkRvZpzLomHc0uL/EbB1h3kMToEhrE52ZTjnUIcoCTwsf2YD9
Wrc3AzOEQI3WdiR2nw45OhsogEmwQkHvCI+8uF+MK6FY6ePVDTPSOizjqBopt8+t
ckKrogd48uPzlI6Ajjn+pgM/UnXuePYNWaaeEku+mDWVYv7zlaWfVfutsGnDsjeM
ogvS8ZC22v1UUhwBfTrk+8SNB2Y3QmqoyUOJl1MRjnLj4VZvZAzHKf76GYm/X7Lv
76AP8tyjnrzIW7uqTRKiYCWWuie+6Iz3SR0nQkT5EcEj+1VwFCwN4177praix4Y9
ElTmqh2Zs9CkIbtocG7lghsKbdsvIuXYrG3TcOTlsQDbzyVIHmJRXqwM5HMjA1Z6
HCuce2oQl8o+43AXbCGScMaSMfqi5NfQpD1+BkmS9gy/warxPVRljmYmJLRhqlia
nHUc+rz6/3VJTRGsl8q4CY5mwK8/RwYYbcDD6YkeXSwX/nD/jmyVm0QWH9VHda6L
Py57Dc1oTF7fm78WiKK66kci2wP0oRNqlAseMDoE2+HSgT4nh0lzeOv5ITrflMfi
EfNUxc41HhFlh800ScJfhF2OntrQ9u44QysJMZfAVC2fFIq51Ela2oG9Rbwbr126
eF5WZhUUW92NekLi6EkknHvRDWpcPsp5umHHIHUzxzr1DyuG4S7YWMXwezrzt0VZ
qt/S1hhj6+x1NtCe2nYL9FchjBTeJEiS6OAvyYDk3kuHbbyeJDG1q1l/U9MOK9GV
wrRfJTf0D0Y1YcoVPQi0pF2d6LQ/Rvjz5IrtbnXibdyk1CGJAu6FrikRD0BVJ+DZ
YK6N7lLXcWq2MGBx4TmwWy5z/9k1nV+mt4H7OVaBT30ShviirYjLTpmhseuA2Tvi
538mBd2QkDgCgDdrc14LQ1a8Ek6afisdLNHO3gHXTqgc9AscalaEuPpe/dvAntA2
lUwnd0XzEY2+qnRqcK+b9tMMe5QeENcf+fVfEgH2WDHAIVZRXzNwSdibItOGXxnt
A1+3GLsmCBJrMZpngxmoA1uOSAkj81QREASm2JIiBqyZUlOWhohcKpL00nIgB5WI
Agep3IPciTKZldTu6/39OUbR3TQO6SNkeHCp29KK7KEH7WlbYv0FLRuyMPxy7J9h
gr8JKOHulMJyslKWBTllHfmoix1oLM61ubc0xinpwazq7P2HOkuS6dqbGwprYgyh
pWH6dNzy/BjCqik4QGev8XjHqKDY+hU8B+g4968QQu25UQhq22NuLWl9f2m9LlTE
W9QfNb9dcCtXcoBqs9W4uC7lsCUIRCmTHrIRvDgdny1GOCEAWjYRi8oUca2qns7N
LwOR/GZezsewlmYhFYUl3YFddmcQH1IpXfiAab1m72fOLTnvdOEv3GgDBUpBZdXl
sovXiclxr/QyhP7D0hdDncKCkZc0aDR2NWcSK1V91hdvoc8UkwXmxz5s/EYyZHXa
03q5PsVe3YdGEfEwH0PmPb+v1lYPT9w5GIVKaiLs3zbIwzG1Rhv0VgrZlOYCEFrv
6PWCoWMWgwBNsY+gXoUvCNhXL5T/JG5x5/vzYV0Rum/3/5emmoj21mH1v3ByVYKy
rN13NYZgxvWGgt3YosFUB8QFUqe3EhWrRAzaCItgR6E6RjDfhubWxnPARBhKay7h
Lyu8dYHCWS+bEDO0GmRsiPkElq5bidEFuUzZhlItlwLWeIL3RQ4bmXuseu8I8WVy
TeTpeJ5yiAB2L2XmJlO/xACoKh1VmO+gW+vo2NHN3rtjRzVXpuiym8s+VrbUe4g5
nq6xvvJyN95W/zIe5PZZ7/b3Q9HeEjTXc+4SRAbEmjNjWbaK3YVcuXfb2nA7WrnM
EYrKr2sYfv0xG2vYA3OlVVYtCG9Kx9hFwkcBObUW7CHlAqJc+r73uivb7gG+qkFT
oE8+HiZCIYcTCl2+WGUqJJt6WIp2A3c1Rpw+Fm3Hkd9/osRB9CaI59n7VQ3h8zkV
L3U+gc+FL4qzSB5RmY/ZT4MMsjF86SKGELb6DBh8wN/dKQ6ycQiHOfg3KTja9O+I
lHszD4d3aE7cIZplevmZMH+urM8ad0+RXlrF++SRkZ2AxWt+tkaeZkEwpSceJFqy
vBrk0igGsR1Y2omFRc/bHiIXPUYNyr2WEhhljMFUs4E2BYJS1PqC6YNfoRb7c9pp
f3a0qbKLi/ZOW1OhnT3lVN2t9MyuxxXE6Lo2hv+t6tRZ7cvXlQIGCwuq5kFPkdsF
5W6I9CwteGkRga2quQmdWOl+wFTZPnW2SJkkeoAG+0LnWCbmdYsVcS/y8LJbh2Ls
OzLPBWWhoSAMv1Lhhks9sUppRH19uo4NxG959TohUpcUDU0LTupiffhjs7By9qIG
wu/vqWKw5aVbsUKLT5czKaFKBBIiv89tchB0bVUbSvHRSIMU4CTCy4OoIgLVHFXb
Ou+4cAeSr6R0kj6ZqDdS9ozYpMKb7jDiDKlC/n5C/mbErXILdhxdZovH8pzFoVjK
z/8uFkTfifbrqK3xbWOvZLz/n42i1aTXXsvkF6o7mqMGxzmyr5EPF4VQYg6ULW9U
JFhPsNA2mrmGd5icDIxcuM2p62y2o3K3Gb5UJAjBtSECT4M5Gl7Y75KAcuDgZa1q
KeVb1c9nksgqwTAqfOBpl6KTKs8DPY9gEchhUCSwDWo+O5hNLDIscgOqiBbLAxLQ
Gm48oty1o0kqeBjwTnVPqqScr+m8FeRv24uLe9hxkE2QC0EMM80U/svQk60s3s7x
Z63C3mikiEXKWEoqM+P4z/9eQ2wqRRWgXZTbf0z+HSo+wWXXUo86VV+N8ph4qPb7
Xcw2occV0SLwckHEt/rbOmp/PCxO9Oyauz2C7iJ/BdDgeTyKDQa93igOfud8Y1an
FmRaVMEXx8cPC0Euy3P5dAerhQue0pmjGY1sQpGjj1vG6rUd3Q3ixPVHEMFhv4dA
Pzc7+Zvc7NAiOfTluENUTkcmDKpXlBHIGP5de2iyqtsZXvARcmfKorowFUH5wgVy
Tet7QG6bcy2sxjvpoyucUI9PPRz4pFivc/gPrAN5ILQGikxqJbnyshSkkAMlpPHQ
odcd3vdC6F+uxZCKFtjUFk87nyohYYdub+z/6vdsip6C/Fm8/MLfjchD+a+jnLCL
lYAJ0MmTFMv2Gmsqk3LYxu/6YdouKblNAs6qlolwZsUYxajXGrcrerMni446E5VP
wegiqIZ84vtGQSp7AY3/EnwQRFzf90/iS/rogHwlT9/83xkTCmfSWlPmmuLzTIFL
v949LjtoCoXz13DUvAD1wBd7DPZOQV+EUH8ysIHKMRQZPW8TBLWq/olVOBIdky4K
3Ms4iYrO5JibKdCUh+7Uc90A0krGxY65dXEoPsgATioff9LbwDNVpAbetKPNkUpf
Xc3PeAiJDUWnvilQXQ0IhFkk53wh2xwnjoAQbPJ6pY+OjCo8b0dFCl0Ei4aSVBGm
I3+F8JKtS2KdtCUXLZjNRRaQ4GcaP2YuPwR8tyJ1bQyz/bEKxsUy9CYdtmNjPmfA
eaWor1gsKbyW/jZi7+GipNFP4pP+NfTgg84jBKqazHCIlfNsWabj4ZxjhrX4x4yS
uHu0l1afPoLvOrMd6/bQqwp+YpvYwHw2J2HgKE7jr7X4dG7bBdVyz90+5+Turq1q
8Z5an5/S+A8V7bR0M7TZE323SEuKLZL98ibCtg+XfBEvRJZ8t5gTPd7tFEd82WTf
tWFoGA6g4EV433ft/Z4xdLmY+QQeP1hbxjs8xIvxbH9G8iD6xad4V3etttL+Y82U
vt3fbTunwBDcKudBX5KdAOSP+DyWVAS3PR+sdgqWyYrxlv4Xr5QtuP/kbaOw9VXj
fmHFF+NpkNeuMxq+NkTGdImZeeAm7N3MVkDqCSlQadoqf+37ntN4FPCDXhObJlGw
yyURcjqlpu82kZvRPAlZCA/wt9U3l3r6Y7lJpj2QBbrgP/GTnZ7mvY5eufTZaSLa
Q50pWCdq0YdxZPbapaEqouiTT09ZadzZcLfYoBC9muTlaR3HJYZlMA7DXHcR/Cb3
pdYr01mcMymvPNIBoEBvJwPPhLfy1VuUsbfDbdI0yCQEWWV4RouZBbG2Z/f8+MP4
jL4YFY8UeJrww670dLdGVvc4kaAAdMh/Bevwhu+4JuZOmeF9GbR1TCW7PjzLGkqF
vf8oUvugrcX/cg7y8FXdRiGwdJQY/NUkUCZYjF33VBXawjk27YwzkTqDDSswsQRe
bEm0ieuThZ5mylcCoTzv7iiC9lselwmPyisWVxiUaC+R51fOnd5Az3JgZgH0EbxL
dCDkoioeSS784iFgYBUDp8kpl5RI16BrUwIlC8Z4Oo/ti73VNebhFg6NmwZoAxvm
n1WpJ9MReRaj/Eai/bT/pm3w729CNsoLL5Solt1ChAPxLJcpS+i1n5GJyWijwaQe
0pdL4SSJvOsHDqLckTECtQBA0jQLDr/odiR9KteKLKMvUbISOmnFO0eF6P0EvgaS
/7SPHcZZDzRvIscC0IW3Gf/aTwGS+uXuAFt1TaaqwAblOS1DGlzEjfHUiwYWF9l5
bsOeSgHXpinZGyDJyxPzJuwruosXgKb1Svo2dsIjVb8aYYozL9SxN5F6vggoXgMG
ZiUd94ysyRPuZyMAZkLvoeAZWITt7zYrtEE/kl7QsEs71NzNfOaHE6gc6GvoV2a+
/S5TVITefGJMlEGoV7UGtxIJ7zgX3nOcXBvluVpH+psy7Q1XH68vcWTQRdELMKtb
+eAiHUZw2ELty6I4UvQHtRIc2vx9C13puqVK9MTmJDoyy/s3qrL1WR8+cGudy9wp
5o85qsmtkcHz3cgsQQ1ZYWDUMDs2UbwU+J5Y5k+QASERlhgaafMD0RHKFJcvRg89
+jgebvwDRuwwN3F3E6tvYSTfa34Cb1d6mS+QlIIRHL7tTDC+qrLfaPrQi1XzoKoV
z01RQp8dGolKyyDKLIAJF7a3gXhhpq1sMOPz0EteFBJIPIqd1e6gZXzGG5kPDHS5
nxoqvw3cUHOQiy4d/9e2POUWDz8F2Y+aBPC+mLs0MSFVBqlXU1YVSGaEFmTsJ1XF
9wQH28rUmqLDxkavOOlZDdG1Ih8I8eJUGSnNLKtlZI5UBhvYWnNxH8alAYu1EEj/
nt257kpbPLoIDqeETWhEhzVEcqNk/qNZy2h30siFiydn8bqbTB54yty2UFPY1Zgl
zEKye505SAMZsePDX6ntG8YHka6pKch5GnrGvIwW73iszOtW31E7ap6RZKbgFdy6
hM+T49u6mK6rCj0DXSQ5N+OzHyQhXJEnuB3UjDfriKUG3FfwEo5Ej7htwk24peLr
s3sK1IKEZRW+NJcv3XC8J4SGJVvs/5CjNOu+S+vM9hqHWIK2N6ygtwSlByHsm+J4
cswz2/hXRBTB4Jo1ZPU40EfRWdODaFHgYwb954D10qL9HU8q1QIEpJX+Zx462XOU
xDxHv/07dyni+gIM7NIkbBcgPLLOVLZeBLbs99ArOkW8PMPeTxTyPCttYuqG1grk
pHt/RoCbsOWLBEHZxHwaeKTuNmyRjDPmgL82K+8+g6DJTqqJ7u1cboxTKmR9vgA9
Y7RdlUpRKDtf9k53hPL2na2oVJ2UDbMiQooHeXxHpKicDVU4XCieVI+vGZmftyhK
0o1NNjgFZDAm/epTQ6/3Kc1wWFonlndg/08mLGco19N9XIPaLtUV4/Tt+gb+OdFe
JMkBoehIOUGLcjEYN362DZEWxPfF1Pl7MUQt7oejDyvcyKuPv7L4RuQUMrUV8vtO
M/NUPDlPduQSs9Ksx+DSKVDGuvmcrsnZE7qoGGsF8pZSfT1Cvo98pexprwUOwZFg
nAs+IZnXkextSi6M/xw3ykHqE7aUZKJlYwiLeuT6Ba9WYMQLVXmGl9KwIr0atwJP
OITvLy0KTWOIoBxc/YK7arwLdx8D9+18uxIxF5/cQeA1Xfy/pMj9VvNdYSs2rrRh
MpM4S3wb+FhLZpoWUGJD6ZBd2Y00s5zbWwoUKwGcAyOsGr2LyT0pIlIUrHBlzKzi
WVKKzL1bArTmTHuOGv8HqLM7YrmsQ8uySwdzmyhUIRLskXjosR5k8NkyZKnCIDTA
tW4TgEzrIJ+GIYUvHYhFiCMaZgcjAT/ey3IODOCduaWsa+roG8b4IEmVG2CCyZza
NaYB1Ax7Ed2M6Bm202Dp2BSFq9rei0+ahuaKXRL88jpIAKL7Pim+noCl5HDkoj55
ky5UbT8Snz/N/fU8vr41/D6TuxEdxzAmskTcBdPkWI96tug1Tiv4Ms8FxA2j1g0e
ZTly7VOoVK15veqSbd6RXAyKyTyjaHSasyd1k3XIe2NRp6m7CerKowj6bADyXA5x
WL3KF7Dqmab/ETUE6A7KI7ii5d10RbmZKMrXfiMe6dcI9u0MEVcRX8XKUrw9TqDL
CPPnTfbChb83oE7DaKxRhXohYwU1Xvctul8765bE8Ate9tQ2NoYiTuqcaxHYWEJU
8cESl+dFGmOu2WYmy+JMl0ZuoFNfuIvolUmwdVzgxjERjGy8kA3cGUFVIY73XkiS
M8HTUOxEhNLB1V1sule3Th0hSu29mcaJsIFdDzHvFm2WpUhUmeFQJjXrmzS0RpoL
2nUi07Iot8hZmzChZac79d5WNiqKLWBAkGFFDnwHqNrGWdrQXBN4UJvVYw6hkxqj
LPI8fialMfu9gcqaiFKWembluCo2pndNOgOu3J8nV13M0M1r395mWxA4xKoQ/yNT
RCnVbYOSPmpD/r+BQjKluo5D5lxKR6AfGyB2rzKYBb7VZRHIYWk9WR1jqCkUjcFM
W1Q67hfWncQmwx+ozqDRaeJLmqJk/Kso4JhasE0DwOYfaKidJ2EeChg8i8fmbrbW
oAX2oLlKktFViH+veoQ5TahDMq4dK9lIRKQvxlIKNwNTy3R5xghD+fZAc+3CkSx0
ivgeYMEQxAWLLW12/5tk4+k5aSiNPXyIBsME4oGczTsMWWqUIOCWnr9K0FNnVrza
6Iyk5nBtSu8+iNWnpKbpyinkGL+QfAOBpbJGyk50nDOBbgq5Rxc9W2e8Ibvf7ObK
XklBhlss7VqGDYdnMd94kt4M1/+kLgGSjv45Pib7dFeYzGKTvtp1MLUVGpMya4Sa
MxU+DjbNhaQOHEoIu7n12zV6nkSsSlzhliByCeSEPd/AQtjIInjqjRz5e7DlG/v3
rf933lyMjHnjAubvnyFrqnWQ5wQZezqPu3lGKkkpN8hw5fii58M0kdTwLBw5I1FS
wil3CjJSdXQ+k5QgD2rPqlZYjLhFGaWrEBYNohIQZS4gbQSOytbKMETMDSupvKAY
YDUiM031XePYtRLxkbdeIdAcVcP+wqNBIK4EhRk1jhuBH4HCLWxIGhf5AVGOdvop
v4asor7FvlkTnPeUoUPx5SuQ3MjhG5Bdt2Y5btrF9lRZlqswpQWgx42mDtRU0TT5
40Hxiz7ICy8FX4Hhkrz5PAAitcvVluMzcpXOknpxRw+H7vRy4IwRv2E335kFwyk/
5cRMfNQwVc1B6tMHXMCM5Et/JN7JrVSzi5b3L8OJN1Q3K4CaMRWGL6RnFEQshnA7
OHFEtOlQR1rYfgL/E4Nmge9ohkNQ0EaBUJfMSC2Fh2aWyoG45SKnCq143JtojH5N
C2jk1qkUygJ/5zHGlZymuvrh/MFZjenwj3OaSwJbbWsuwFyLP1OGmu0rqGRRsD4G
RyGfZGR7PZNWBOnzmku1pwXnYl/26PFzUG8qgia/2cOvNHArIaGao864gjJ0P+M5
gIsJrZaz9jLe52LshX8lP+LFeNaCznmX9uNp1foyvU8Iz8z/lUnFfvdgyobQfAOJ
UQQOZs3l5yky+nKVi0aW32aNecwSHMkUEDri1PeroO7ygnDR65a1WaGGrZa63JRd
PTU8vPKZ3QnPIHUeKUwBuwvyMgI9NhhRy4ev6dBrKea/1Nfqd+cJRqn4f1AsX0ci
/PWL1eBQOL54yTGWkyAvA3kUHlGZW/mFDJcZXlI2KMmklUCgFks/0QywuU85ydUz
jizSdopOrvfacJ5bXnBR+SH6G1QoN2MJTau+Vjul45z6JrzXWkvKdhWS5WLP94Ts
BgKnXcxkeYh8fUKwDKRpXo+nCLVqs9XlzyUEQY8Ac5HG+xo+o1tqCbSrewhQIbec
dwqrWwY2E8BZyOQ2xPXjB/srt8b7qHIFDBDC7T7U1JY0T4AyGew1808SH1+cFOe6
XtZU2djwz4j+Mv1DGE1/CzUgyBWnkB7o7URlhel5kZw9D3nT/5mOH/K7iydG/hOi
cLXNp965WL8VGlY6T/i/7nqxTpov2rbhtSPsUrldHbaE+X++VALuC8ipJYu+XX5o
QyepMx3+Ar2CFi2RNKamilVpnhz8YYD37zI74d+o58+8s8dRertZMmIHBzsoi4YX
UtVBS8ry46NrB+6Z/+HATqVtWCp8m0WezLyP/e7P9exlwx17lXsSBvRFG1lnEEnB
+GBoe51iZB5oP+ze1IHwS4GSKOaAYAZ5nHLGicoI8sPxN5KsprIyr5z7e1XOqq0b
IjNtDI9lPGjOwJT/nNHxrEgmFMz5u/4mkr0QFr91bR6UPh8e4x0lg037tIUqv81R
/OKSVQiyU8iuRrW4xHJ4b7gQvWHNc6OF7psYGnBPc7r+GKuLxhjaHhbsINem2ykE
KMwaTcPhXwJowBoeD3yWq9D6anCLruGNdpqiMDXNxq8pWufTN5terRDPy61o9Rwm
iYtZxSL+rGeH/u5dxhZiNLky08eGaKJCtJRiH2CzvhcosBEMpP7GcvL80eLjMNZv
KbM7IhylTTJYoyOQgUaVKdurjG+L/noLXmwf/if/gzWb2Kmou12oATgYDlAx32Y3
XZOC73HvHpRQSYbKAGCn4EOSWzhn/pxVtkvrE0zk5S1RvdDX13l8j10JxJMQc0yi
A/FZZ75E0dxwEKfhZLa4k63DeQ3IuT7KlVAWaOhaHw+JRxrP0P+/7NJYUkz5ZKu7
M4AeP67PF4tXpNEO+OEiMS1/02JtkkH+lAIN1/70gDTLXXgyJTfKaQHiXM/9OK4J
yZztCR2Ywes6F5y0vUZlHM453zwaHMOuDwTNrWyiwes7qhlgLZWrh6cBcL5qIPIf
+T7hDIS+m/berMgo43vhrdcvFwXd2JB3YT6cJXrOk6yGgkqmwr+80vED9YxKTjRu
SYA0QhNofDT4VOcX4p1zZJLEbtYl6gP/+Lk2Xw3dijO1qAzgx/LLLtEaePegYt1Z
1LFEhf+neG8AGpTts9X+oXc1JrWlNJOfJ6FfMVHx/svu4T8hMsC6YghN831Xs/N0
hqkcw+oypjjbOa46vgRK0lyI/5a6mKhe2OzKYap+o5i2do6FaqTFGwDOKvnPNHdI
/1znzG6GONmokqsNhxyG4y/WeN7Sb/0Qm59Mi+I3xv25E3jLuWFbEEspQRhz8M9M
GffOOsC8pRJv5NmO3nOXDKgh58bB6TIHURNjvoez99uk7F+BzqsYbyzFUyVOEuXQ
TxIG6NMsEAL8iXWORYnwNuQiEm9aO4U960gTI0QD3KUcQFlD5B1AMCgdm9ENhAC5
6UQSMIYy9onLxGR9psmZ2attqPF7FJqFumrLUmeU88ycJ0NMBK3wPhccHFm0D9Hm
PZVHSnPLtwO9m323eqPb2mvpEyCe6Hwi6GUqIo2DGknOfZHb5L3NWipdAXSYtT03
GPfYKscD0OiAWfaSZcT7lcR4X8+PrXZtcpAf1t5AG0kGzHX1W6lG0B/+3TWZV+gC
FWNGolaRC7s/kRUEXA4B19D2dCqI1UU9tWXRk0ZUlWvaD+DMbuIX2BxJC3w2kxa6
uqwAOB0UBqIOnLOLApm4oJxuqyQeF69UG0i7xaAU1wNBft93x7XXl9FCezdPUoK+
Spn6YlLZ89N6+ME5CcxkuFN2XFNWACaIPuV60EZ+5MIOL68edZ2ARFpvUmmrzj4k
ma40iEuwzSoeCg0Pg/GISywy9oPT6TLLPyPB2J849Ljsm5AhBspVSUxWgDE8/VVJ
y4G7GIud3PKBfp6QDoNzWGdPkNGfKSkydMK4PvbPrvfBL1RjVwSIpE8dXpXv/2kv
ZGsO4NQvRzC+lpdpvw5W1IMha3lq78sYSrRtZDApE+WEBy0l5BMDy3Nsi+Tq/36U
oRr+cXo394lax/QMW1Z7OTaEo08JPNLZITkxeJNPAeNIeRS0fZf2HExRwumkG6iJ
NGlCRJCCWzdM0BhDIvQKuGEJMGch/0DJhRgPR0IXpEkq3JmIilkqOO4xkeiuppgK
/DHxWUO6+vhR7FhwI8ybRXLKJlVjBggJS/DY1hg8vcsxasq0XiuYB5ObTWjo1sUU
OoaOgPAtoXleMRzh2WsObuM+DgWuauNYYPx0swgZ42F13I79OwSPuSUgQXYlSu9/
l78pYWx9hMatJUeA5wTnzjr8vNIWf9na4MHx7FkMg9gsnFjOtp6KIeiuYwmhVwjl
mEzmKkEX4jOS5pVkmtLTTf6OsV45dINbjvAyoBNPIdrhQTrnT4PWiLFTmhcesn18
pwD7Qn0QEh7oRqzIKoPF3rqX2K1p/pUFyR50QfvF4DX3inh/KzzqYHjLtzqMDdid
UwsNxTf0r1DPoONZD0yWfnFxOw8GhTKrwSM7EmeKu0ctcHq/rgaPqMLXof4aEbV2
jJd8JZNFJObSTJevnXePUUpx6/H8f5itbQbVcJxdg8s+7eOlLu3bFNNqqwJeyPzD
6iZIXiAnBwhVlE6BmCvXqOeke5ZnsKzwQP2oCHpKWFEjK/X0HO933EJjNpfbtAZU
PbyM5tzDKp2IgY5xhVNZdEBewzffiUolAaydTcTNkU4KEPVnEHzHEmnIKYipxYmp
YbiQmDulL211MgHSSWcAM5Td6+KkjhK0uQthKRwbS5KO+KVpImA/Rg1TexZdZBtG
ZwrzwfwNLoEWUHyYCFjmvtXwTun9qAyYEQx7Fp2nkPuAVp74X+bepu/358O93vur
l79dSr1im7BuOx/H3NRMDCTo06PTHfvpV7VFIey5isiLtS7VKaZ7+4bqbyYuQiO8
3FLFcuT6nQbKZfaNSzJtBaW7eVzhRn0zg9rxzA9WSCU1dn/2CX88jF9YKeTj7Ny2
HGxr1rEVNiICQDSmtRTntwM2NkGRUqwD7OF0uxISbSUlUYV1t5OlZcu606Pr1CoQ
mZ2tGyxqkoOJsq+g5zjyzkXfecaqSdYHMUWkx+h3zdAa6J9QfSzxofQWY1nxKzNk
4bAfTE9TX3bFH+S2DACFzIYVwEb1r2L/KI2ADENMpSiQHOj2ySsM4hPwmI1TAElA
uF2ln7+Eed+yDgM6dK7kUvjZO6OeXi3XXiz/qRC+9Ky6q4JOsdWGlxZIpJOAvSCC
3IG7p+0zvSXznnwQl433mbG+5TB97ySG6zJ1bgV6aGqb/nUkWsohdsBwj4T1RBJN
6W/JliS0zvqsMRUqwALPcjsXFnyis0KUypospnzfv9mnCCzwneMgPmafvCbeXyla
41FPezwMu/ezWok7xfgLNbjiJp+uv8f5a/ZHCUzdXVT5AdDoDswMDHSE8F1se/PY
ThHpZHJbFNZpafVGbl38Lo8gDjBF/dJ11jjnHhIODeDMrzuFBmE4xKXKmIxL8PEB
U+kE/yT90HOVl1TdAjCqBrbNj+hj30r5BKqmxdAYGP4wZAEuFonZzdMk+taL2cBn
KtnSEPzo4Gsrl8yVMYGThIX2voaPEM23XJuqBpm9Y/0dQ0wj5SQR4Y0kyDPDbxUT
HQ8vzJlms7paSwHg7oKRJ8BVFAYPteB/xYLg8NHfA3/aMQu+fhW0CL2GA8gWWQf2
Xyj38btxKsse29yz8NRdsy6Vqii5ZsU57rw7EDRzSumiagX90RMbpNTjcdyg/yt0
W0lBTvp08r+fO+fV9nmNVwSpha7VX7rOjGYpGL60bWJuh3j8K8RkDPZkvkmAS2Kb
wXtPW4RsdrsJZWZmRF+53ztmou6psriJyJOmsoXRn7qu9nVIkySo1rX4agAx1vK3
e/N1rCxknxkIo5RbS9JAzyGhz7GnvHulEguFJHdcv4XM5GsCpy8lthlO3bQWzBlK
zhgqx+5X0UwkESJxEfezzVgyZ3gbuNyRbIe9U7Ngr/pjxGS29OYQq7t7p0Op6ElU
uZlDwB6jp4BlF4kniuHuZEiDi+i+WvYRx1k6LA4Yhie8HISoN8/i8/quwB7A1aQr
9y3OU7Rj8vRtvXjZ8lz/F/ID3QGp02vUzTDhvaW/tuxHCPSryogQAN0UTmBNJlQ/
ngu7arkWXIBt0Db8dyHN0hno2nCTFSUfRapHl4MFB8qfzIiJAAz3C4SeumcBw1pB
YI937qZjx2wW9kN9bYt7TdbpGZnaoJwug+oYNQ1A+elGVZFHwdBpn/NUsu7lcZGL
TFLRVY27BOOOL3IZk9FZ+mOPVRQOKIidU6FOq8166/j8zhh4pTdglzNyNgZeQ4pq
2lBNg4taMiyDLuLjPhWJeXmbZ2WYWqvOaOi8ontmHA0mYGNhVsFxsX1aRSzJrl2Y
M/3xj8/F865p7AKk8281A/lmIYInOm5svY7/P4oWcZZKxJBAqLfwJunWBwC9fx8O
URqrXMCFRw5bxU/qxSsKDOW6NlfpcEOcxi0GoVxwfib9Ah9dYb1wW22xQJErBmmF
pioQp6FOXb4xXaiSVOp28epKO0B0dkHxEeI9et7vk4gtDNzhIEKAUCIe2IKLvL4d
eJPKOiyUmmYmk8XtlK5JSPmCdPowcPA7Urbpn5BKO4mFm72mAxzq7XnVuy3q48g2
P7EnTaGEWDibt/U9dhl2eV0VHpXg1+KKBE47n2SB1HLC5TXJMQh4zuj8e/cqjofx
h23sxTJtF86cek9nI7SHI9ZLT2ofJRFbzURi5+HbB8UZK3FminV8tIam4iq/+dLJ
UExGtV8AaQeHlEYCIfm0gfvzMr6F89gcK1x/YucVycAY3UVvn4LWk9xurhqx37AI
YKIpLmngIaP5sSXHnFtEBmX/Nz9ZxEjsJPwBpCR3QI0fUV0gbuPFjZfLE7GoIXyo
1fJGeZCbymrCntZQv8tg5lgZkh6sbu+XINyLYvoTDp4SVExjE3/exkVT+94M3vPZ
OQA32Cm+XQa818VxDHDQ87ssfn0WNwjhtnjkHrh7BSQpWK1HCfzSXxzElTCHQScj
UuZrUMFd8xOH0YYcBT2rdca8OFIsJGXkPwLHWHiZW8i1fwWo6P96j0DkNez+3Zq6
Wx9NIgk8yC+jMkLAZ1FpDUTvPU2nVnSTncBwDZsFIs1ByJgB9TOw71IhFYd+QE3U
OVbpmSAgRaByV18+2w9yQvUm0EK6CBiwSG4mfZHKVk0PmJKG9s9wqxt8r0KQzJka
N92Als56iWSKhA7uH2ilaTWqWMBQEfST5BIrvACiZPzqA/hj1Mv0z7rNyZhXYS5K
03SLzpAAj3lIEFFoJXiZjoKtfcQrzMEtzju4SvVSK1dcH3/eZoH0iaNy+a5hBYlu
98zgk0e6mMQaCiM72dm2M7KKhZ9sbbzvczsDwoinidxqTYV1d4EcMtlFc8b7RVag
QhlBVau+AxNjTwOOym/F/5inRKUSDtT3ZLNnFaRRTiSHRjBpSgYAx6YF/HrGRX4P
raWlNCr8y8swJgXHKvyaGj5pZRzJBbtB2pHGRqc7ol6Qc5JHb6d9iCEk81IkskGE
m11Y7vANqLu98t+oBREcjV3ShK50ZdlQUPZp6HTIxA4Ia85FdDAfv3Lke06i79QK
2xOEDxeS7p650unzDAX0nK50RdmW26WqIDF5S6++VOxNpdmk7+T0A7iImxMVjFr6
hOvuGOuMbWBplzkjbDwbAjRHDPiDX5J89ujBuyjXOueCNYUke4rXnD7SvTXyxH6X
XLkyQhKH4jtJWYEzV02wpQ+m0T59Uh8XrKzMvRWcZIiRZx0kPikxSuI0Vb8gDGib
uvmXnmBxpfuCN8vznRbOkh3yEqAG6uUd+o1Jce0ZZFpCBF6+hqv1Rkb9UiXQX//A
yi3ULCPlZhKCdg/9CQLNgeJW+PlslGqFRpxEotQqF1Vl3b9ezpPwRFqSfhW95YTZ
F8XoVuZLqO7EnZRdVK7tPMdoXjPFAtqhgC9hgWoeuW5cPQpRjt+bcnnZZSbF2Glp
4ry0bnXW57YD8Hjja0xIIhaY2OTA3CJG/E1bnO9yUIjuqcwVRR7yQ4SvQY1kL0e+
BaysqQrT9T1ImCbqJ6HDIRE6DgTnFqDs5ki1tE9ohR1IZwehtny54P1cRNFUrY3G
kyPw0v4OCWVIrniv/OGWszft8fMU702fq6bQIYsHryDNGOQ/jsmdWxUvs/lIk+mE
WrMcR5BJf1CS1tjTltl1mQeJR7ug1SaAHqf+vexqCxGSKZHE2Bldk4RXv6IAeqYi
3/og3xyBA+cGYE1ZmLeqUVKNJ30UW2YpDukdkgMYl6WKqJi6EHkcu6hmBG5ivvWS
cLVTpEVbw0GNt/bSgnHIie4oQVUN9tzfYByi4nOkq8//hIfmCbzul4qisgzD9dmy
TndDuJy/FcyDd7SEd+WDjkw6w6H2BZh1yJ331kkU+1BJiixywFP4VeVOzkDA8nf+
pJ60btZ1GZMpnB080r3w78cgvmFhcMSSaHTQGCak9rfL1PUUuEshp+r4/jelDLYa
QpoQvX2O6nVy2e3UGai57GUkn9bCj6pvF8ekVDlBBrtpmPxhBJ+pDfIapMPyChmi
EMnZo1srwWXYLjdbsZdfT0dH6StGAZJAVrEOk/lK8YMHl4W+sGKGazgRdHM7W3xn
/6VJuhStrhWPYuilVNsWVyg8n7p++79fHw27KgSRNLKIPzfi6tPXrN4VpGU52OSP
SYkPfibE96cvQAnEaynP37JY6Guty5YSpwUO6VzoGuE/P0uX5Obzgzkz/vf4Va7d
EjIu81WOyTtx7x+ugbZRuxZ2kWNclcPh45LA75AOomIiv7RCSSuWs+Xc7JFPxtYd
khtdGfclB6MNjpqceKsObK+3Ws21GcN7hZ7iWouIWK5MPq2EuMMMaWVoD9HrbhHD
wrbLYag8qL7EFqVq5uY4alNzxkggWPSAWSwUmrfoP1ffTGvC5IJqerqyglUnK7SY
aJJj2n6qgNTijCymD+N8GXc4pdWl9Q3bbUyFCboeHKa4lPA+Su7IkRLrgykqKqN5
E/goOASSMrDZk3ac5+Ni4r51Ydw8A9caMqAfiw0LrWhiC9RjrluF8G+KQH52xBXr
4vO2kA0sTTz+Eg1T9HXj0FAeqCq4k7m/SofcQ4+KCLee1Zmudqx9VgfBRRLnssoh
zXMa9LguWMR3LVKfRmXnTwBNMJXKR+7P6twmJDHBORmyW0YIWE84C+2Sq7vaXSDr
vMdkVDGAf8l4/kVZu2nJT0CUtWSwe86G+tuCTn0BbOseBhr8WZ6L/rU2S6wgEi8h
oSVrYKSwEvrgjqNWNUjyMTpWLBT8l56Kb5FZ4ol2atMnbavs+cj7y6Zuz3riX2YG
RnaJ1IPqzo8Dl5Wf9qlmgyQ4zMK6AShixQ5SXOEWdW3ScPo5xpSDz73Uw6nZn8NI
Fmr9QE+kOyGh1wOPYD/xb+kHgdrWQKWUVh/1NwXi1K8cwXT4hEw24gI/dmKLobh9
NrYeGzUQNjq7zidfOfo+/jdvvv9nSJ7k5awlbaRYW3/dSdCFTZnUNBNsqyqJEYZn
J1scnQl9h6gFq31qWjbbUHUQitiL2d/1U4agJLhwDYUiEQii4ZWGwvcu/RFj3Ruq
zGy6QvaeFZPBaSbRwVnfq9pOPSgcN+P7W2Tg+v6zjV1aHk9omOnE5AKgYeh+MiI9
Dg1pz8rdHrqXNBywi3d+635kSBbe52e2iAF0n1L2KAymAGyKqHmQjc9sCXZY+l0o
477LmmLv5lbWv8z5KBF018ye3F0Dr37vNYs2F6k8Jo9disTchNq8ZwdUKc1zKaQf
yLt1GfruaB/K+vuIIblflhqMJTSN/P25We/R/Nmm4M19kb0BEZMGMhTmOecqbKZE
RSmWfOmUa5qLyQy1AAlLenAOoGn44Nettz61R2RVRv0U3lOAprD5RBkkCmpOLcmp
+EtOsW1LnfnBBUcYaRHfiqbLBWoVf3yW1NDaZWfvrDKoml4bK1My+ifw4zP5feIN
1N4r+utbAtsQ5q4B/zj/28Ncacpvv5/lj2txsvkVe3fXXIsgZYb4YyQiZitThMYa
B17LWyGB5bc4sAUv4x2z3gymZHUhhM1yj0W6R0CVdXhsO3x3w7/QaP7UWrFBWnZg
7e1ayTl18nYeCYcDlhU0wqvxyLMX/7kWDzLmY77liM1oDNLBrCf3kG/+fFlUQnVN
rkNrHKaWkkK19ZtOVpgFmzIFzlc2xeaAIRRVuzE6txQTZgmQvudcIrFCEe+ypd5G
H9ZdmU7pjveDtEtvm9qjyExxAeTIQ9bIkYi4T6I3giZu71YqCjXWzgVCcSB7msjc
BT0GqfleYzK3Q16qn7YQvI/oO7byu8IU2+6kmHpFxi2SXd9/Vfpy+bvMSAQvp8j4
e+/cZfFteXgD9uzVqmVOo2NNQJEqhnl5vmtrcV5JFbr0Aqss+YU/Mvxe1uGTNru5
xSYDEW9btwhxdDrNsDvh4eBNTlspQMl4tpDk2n5KY80lnd8BywagFYbINiltlqAF
rI5vzSMBH+LXAj994lEN1w7pnjD59OaDRVuE/OS1YZfj216zxZxGn2qwYerH6bCM
GnDm/vpUaRY9ChXRQmtd8b9QKl0Z/eWnz5BVnVtNuxRwg8L3OysB1oZyMDWDRlOi
dZ2cI+hkwanR7fP+vlxN9IovvcsDM/qnAlKgY+WwLfyyIaeXrE1YOpbyGdvjnHWE
EePOkmQLXyondOUdnR5rjSJF8f7+buGLHr8QqQSTYxwbT6QPXqDm8qDxLRmS0TbB
5u2PAEBCRfq3dqVR/EQSGCQmOxT9XtVY+F/lWaDZ+kT2kTVFZwAyAVjkqhS/vexY
X6+n6QgyFP+pSjJfc3m0NDR1JUuBes6c/yZ7J0mCTeFIQ0a3AGs7JNCj+Yz226I5
x6UhmLYIMd1r6En7cmqlWxBcpiMaeIm++0/ItE0UY/1S9YmKC9dteu3jSFCVn2lx
wOU13sbIXBRKG/x68sOaxFDLg2pdSCYnMs8HKPGVAi7CDfs86YRD0P9gmPJmXgtD
ePCm87bQl2EuRQ7MQ0fPGCrjrX6uxFtsL0PUfhXnAyO3yxdi2M27fU05+wVgaX+n
3lBf/6BOVwDZ61s0Y0CAbEZGdxBz45COWR8VuNqVD11Nelm4Zh0ezMJAs4y76wcJ
+1vsTLikvmRi7ybyRpNASVIQaCjldSpFDST9CYBZZpB+eSJjGHuBhk1hADzBmr1l
UgcIlmhmQ7N06iLJ2rhKH5ibJQgvL3jAMYpuJkS7lYhR0KrKzr3Q2dlfRAeDfcaO
9Qk3PPbFk6dfpZ+chkUDRfg7dhNiDo203lxZgEMXNOkws1i9LIjP9UxgnaITwTUx
c9R6//fEbyMyoR5Fhv4D30miGpVLPvM4tefYOvEYoBVbmMADtrkXEClmfeXfHppF
UXxZeCcgzgEylTn+AzC6hL7Su8jy0t3OqWjuqaUXMZdo3pq7786Ybs/PRPhdgr1o
SHCPVMa7aXyRnClfsLWodF/QWUatvqZhC++XYp75j8aL0RSgkwphTj5LOD85z6dr
8UKryabYxkvY0urSQq0YjPG7JxtJQpzdaCuR2ZaUPTWPI7Phz90gW8mA5YtJBoB/
+fxyw+OnO9n3p/rIBHHeJOMTAc49am9SQK9WEsygBM0YL84MocU+jvfaVmbgNhDA
mTqzlWg5dkOdwJs3tgXwtR0HoWdK34VnVxj60vEVJtrMDAnnvMvEwSALFKCKGCAJ
Jj0pHTIebRXHnQP6HdRhROxmLqVJUV3D5S1IxBadC8TV5J4LzrFj16eVgx22EGBu
GUZq3tYAVijck+RW2e3slImCkCw4T8kw3PgU2QhxhIvWZ4tRM64isrGkyVRfBnmZ
QNsWfYlaTFWMzeErCxn74pViMSPHHvWU8sUTEalHtD+1fDuIaDC7gWVKvtvwbfmt
gAADOX05+vTGMtvuqyNSRMt8Bi1TT0pD4Uc+5g45wqDaf5nUo9AcFBnkplO4cX/e
pNC6Q2pozMPFFzaAMpfCIVvHRi/0q6JQvbCmTtZpv8nusvXhBSAkBUcuIt9jZeLH
Iu2P1uACmney6lpTRAXbMPjXQc804HLh3Hu1ytvEk9DBLX1pIx3C16WBUk3p+2XJ
+cmYtWWr+A+wnbcojXFCwmKxxuG8fffq0zyJc70f4+URNQ4v+7fMXXK3d1aKfENu
SO399xYKS6ef49qmxrJdL+sshYY0/bVPKAHQ+r+2aYtOIP0BB32bDzdXGjIXc0AD
kMDJliqtx8ABycxn7uxtq+V3yvXnRO5TWcy93z3njUAoK/uYA2B3mLx4BQllsuH/
vpOplMjOMzudgzpPYC0wb4G3uOLWt9dEOJ8ePACRupLmMx+zDkjFdkh6EeITa4TE
FCtzOnrhTj1Gr8x49kcuxdpHIdJvl9gYZCrt7nU2CZOPPhrASMIsKK88d3tpR35E
yGhQnCwmGoiSvkEavqeIog0rKg+NRQ6bPaDMIrowYv7tYQNLwPyG0shL7wMCdVLm
2f//gjBhobQm3K8qkkJrXX+Tz2L4XpcFe6CWGwQdM+cShzpHH+xjbwnGYMLX1hVV
JUzdysOfM9nPy3PnLsytakA1Q8B7UfpTtYqKGoiUN9f0/CMxyjQwx/3eZM1DH7hS
nWEFkq05dh/J8faKwkCQt7rWumwDAQ1ZZfZPTpuw5JFIRZFj22mSrPD+eSN/ehH/
d9wFG/h842p/frY+8W06Ujynfuugwsejn/z7B8Uo8HfRmZcLUYjpQc41Pob+X0WI
S6nt24jAT8jZeUecEClTt/w2rlIakQ5+uzUq5cOL1r+TLK3gcM4I8KdZfef96rqU
hRIBUmRPe6u7Z/cTZ0vGXTGuQ2vbWrVgHw1pMHWQzwVCbYW/yofx4ocHZI+i1VHh
pK3v5bjFsKfuo47QLrPzla8MqlKRlL+5yFCWnCz0UV9LxaQDk3mv/Dz8RZ7tDtj0
chdgGebXq9MMsdAzp8Ba5Dhazlv/XfsqkRdswnVLUFfairgGEpW2CTo4DkMCUMzG
OxN3wzJCQVLykE2xgecUK/NTvkrRflBYH8JMX8Zc6R9Cn0Og+/RQImlz6hdiBedd
1p1rRmHkFCqzVXbJHmCiqty6HwaPGZjMtvtHsO+n0mQ+frSA2YPQXmbchYbJLM87
lk11TJAX6/5qm16U/Ec7XFhKSi882N3zwcEkfExd/z+niheyIooV6ZJ869MiCah2
1jncbmGwxNUBhPXujGYGtN2IcPafu0JIxOnBrGBK5WfxTG4cO09rHVSMU16bbtlr
HBhViHdYyN+1hjk3Ak/+WXKeXFqcGJLom59y/xN43YtCjXO5h/Qi2PvEaaLPJR6e
dohXJWLwAA8aDnMYVxSed0mao2jjeL8S2WJcCgd05loUhA9vMZJDkBqO0ha8IXAt
mD9lPrVm4fG2mypKphRGpDXvxtyxKRXuhzjZ9p9BSdjdC8pj1LAdStMphfRkvLij
O/jnHE+I2STKImsoqo0Q1oBc0nLOcm5r0zeTMlvcz2Gb2AH0bm+oGdEuplbpD/MH
l3eML8ly998HTBq043KWNGIOyA49091+hXuQ5sxIjWkoTrcSMsy6KzSr9MM90gKe
wXqEKgznmgXyEXCUfIjvstUm96CD5N2K2Kp8MEZNcl9SqdUudjfPrD0Z7j0n9DEH
EUZci9pQKSB1r+7bgaCfTC/yLk+vmueBfGV+rc/tBeASyttcVN/Jub+a/caDhUNY
g5Kvm+qozShWi60jinBWsrZZt89hbtW9V5iLMcYuAhlZjHzL8c7c7Z0J19Hzm68V
Og7tOf2OBIaW8dqYyz/fyW4xyz/C4xs7M0HC4P3HHd7Si5VqsydDIazsAQUP+Z7w
Dukv0+j43Ps79IBwGSqJGQ3pX/1IRhV7K6nw5XSmAXVQvhz0CvI9JFxwyMCOygpm
JIRUhcsHsyux9uARLuJ08wIXIPy8uhACCFmeLitkEBt6n05gTguVlM5Qdb4gDDp+
QH7eyeh2VZU6i+9AuEFXJ9w4gxrqLETmv6NQuCANdcvocmCAOhKlC2wXgN41Q1XG
BHAIxt/Vw4C7yt2c6TEo8ISlKw6RDzuiPfWYI/i4kzzfh16NAJVTSK/9WVETn1No
dVaEvai9IASY9v5KLj/F4rkbxFByMtJzV3/nQUyALGkBrMU3T9kMMmiy6buY9jxe
a/oKjOlntiR52X7QqwpxBMZovGmfzw7EMF0Rea4wQGlQfNMfPB0HWOwYksGcVeHl
a1TqYBvjtUbb83+Gz9AaA7K4+iBjn04cHBMJf2WK30qSLoBE1RSk5F4571B/YO8G
JUWTAg0/yephsYIBLUU7kWbpXN0q72kwcGSLi5KVPX6knvg6UciHM6OW00GNtSHQ
pLeZZ0Ye5Sh5Z2MJMmUAPY+ywGVTezhERK453i5enz/FT5zJCgEUbLA7p3/ZMRoJ
+XXm3AxPSrb2l7CoxN28P0j3igPhjE2/ppko1GLSNjlsIV5h1u3H9xJmB71dTH9n
iBzlhEV1hisCXYdMYa08Qz0itPBOY5Crv7C3q7PXsGt8UUDL1jksi5qr9hF3GVQB
4mxLk/1ukpLk+7aUF3T9jyIbgD+EJQKGs4XPEpjRRriHlIoFztQoDgwhkVWnoczc
SQ008VBSBX9wsHvY1XcG8u8XaduOczCKverYn1oC72/c8EhYD4+THHWOIG7V+Pdr
k9cilfz/ooA3PcfQnu7agGNhSIr1cD0VppTkc/VUfA+OBGzUInJKeS8mAajqFOAe
ofXHv0klFCvk0a0sKhuCMThUarQWfh/edxAW5EW+uiOsrUHy4z8rKy29iDpIAzpv
aSTGSnueTV6n6BjkoNwqYwlFm50KOf6+PBb827KXTtsEeLCPY+FEPQrcYwj25XhQ
LqV//UFPd7YVdUZL/URflbEreIqUXgsZddnRB8/6PlS57hH1/UsRrPnatb7u//40
K7jrwPmRNchWhmOEjME6eVoNnMMl1IDzNupQk79QbmETO+la0Bv5/qKpibwaNh/b
9G/LySB6wONIAWKnfh3SAHbxnV85wYBbVMr6eHE/YZqswkxlOMY9GjWoi0+OrtKV
+EnkizPxxniCpI0bgsdM27EchbYj4uNOUNT5Q+j9CBYoTf+MpWWk2nj1rw8Rdp+5
j5N3QZaEkDrSfRtheHWm0Sr1+dG6zVezjy4/2iuv0caPh3Ksr1n8Z6wrA5sA6khf
fjNHd7dhPdYQEQgwscxuiFjihmQdyorPvv1VwrwIPCHEI/GJip9W9K5SkXOXp9VH
zKAIEPSajZdQ6RqsbI6YWdd8d1FtiuksQ1P+Azh49KWnJurglpSFKDTi88E6jyFS
3SQcOe3FZYfCBMjVdnaOwrf3RhjwEAGFAym/wgwnAjSIPgfSLFN4747F5UGow5G9
1gqiEpT6ZnGA6xCcHn4/oM0hbNCH/l1GuToIzfQhhKjVTA8TsFteIN49Z+HVsXZe
6frvXjAeDt2XeAhEgd/oozdka7RVSGnokP83oKLtgAZGsEq+BVmqLQ1IQ8BBNaTf
OZIzrCQYlWBWAv+onzuHD54eNxO/RsNl6f66037L2HgUrfIJyOBVJ5ofbmoNOUYG
knHGMopGfjzFfeS3aETV420VvwG+sJQO0g3/Lh9YNQrMVq16wNqgMv+CE+ZaD+4a
evwtBKH2CHhf1/DwphH3mEKSgaIkJc4Z9RpiLw10gwjHpjSvIFVHjzBd+eNBkZvS
X/Dg8IhelCuZWvYIxzYIQQCZcub1OYnnWxEvqGcZFBsW0Tkx72Da6OzXltBzE2dQ
4gNDoQaTtkZNECk2E0LHiqwQeOiIA4iqQZyhpaA4MzdNiESMcOwStb1bfXKGH2YE
ufjmIz85WfyF2qt8AAgR9rWAuTRcKbfrhi67d1TvBIh020rjly7zq0HCWatOcThc
J989DbeFj+Q2TPbP6z6H6pVM50C9JzELfrNuQimehCkvgVcaCvC7//TM42rhc/Zp
ymp+vD7ZxgK8M3Ytg9yV2D7xSwI0T4dvyqlVBIuGfBVfZH41UEk/a5bVz8QBR7Yi
45vRvzFhBIyBsR506is1eO5g1dP5qYrHm/TIYRgu49F2RUGDBlPqPoYjtlkTx/+k
wc6wmmZoZb0ZQFcHqBBgAaVn+bMXClazjPNhRBUKN/H5aTjvTSxSOJQxMrKz+1NM
sYekk+J3A4MC1XGh93hgpomgdeadDTzU2TWfsj3V3KXz0AOlkHsTmwpjxdR3xkLv
PqhUMPM1dkgjwXME3vPG0dA83d+8mVaKoeImf2rHYKnF2xda0Mf4hiTw7ZAtEhLp
KCpdR6rldTQO97/saSB6cb597Uuk0kncskvCxw5h9fjUo+tL8cF9Sqca5LPbLOHy
9/xslqVrH38zr4R4aEXtJSsy7BGQk7sIFkgzOvt4fDU5Cq9GEsEZHfYRfnuxwglS
aRjjOPc7/K/UO7QjgH+AIWiK16zAy/CsT0OEMqqzxwd4yb41pLht+0LBVw5crOa0
1vbNE0XaSSwVs9bqohEPbscg9LsSddpgtgcPHpexLMPsDZvWGcy223y362A22RS/
Z85sGfGQLNxixNThXF2zMT2HPK8VNGeyT3W5h51JvL2KqZ8TOEvy5v6uMh+/qhaP
Oqswag/+dCkqbzDV9b90isaXHJ+NDcw3BH1gIBuP71X4Hc3XRMjnyZOCUjB5sgAI
SIMa6xP6w7yet+BoIr83b9gfxg492cqQ+x9m08xhjpfbMqNfx3TOSpCZYgOwFydl
4zZ9jeGjxuX/C9fWwIfUerzQ6lMcj/SvLmLXBlPj2opL+IPadtwuDijVSmpWX/zL
S79I6KoWppMbGo6IWk0xLtu/AASruRo27N3SZfataMDkrHV9PPGgZk4P+fErJU5q
egJmuqNbUvEz31ZyNb6IoNVoaD7BhyM0a/IVXWUFkDrCY42sKWXZfEGCA8DYex9d
skhKoHeUR49cITkMNxvcVDuOO9mgVCJHqSwVrccoWSaJD5+LLM96JovBNVAGbV0z
yW0vAHfG0JY1KsEIeXktbDw+RRQIlh2Xbt1eqUdDJu2I0kU4ZznTZQQ6IEI/Gj6j
smG6JTF74GtrLsjQrPBLhDru2aMzXpOHpDs/ZM7ZXTtSKpURjwklzL9E5u7l0/j/
sgUKt/xbPy0BVYLJPhx7ppMaXwU43XBcpkr+4Uj3g8kaWwZDSKCULIiRjxdGjdjX
nF95xBzJgBEAkO8T8md0D7H5RaUhbfa1n9MZmtoJoH9InzSIGCtRbxcJJv/EPUJ4
OfI2lhn6yGn9ds3rZRkntffMsTLSQVPvEiR60KMXa3h+vNq0bAeUZLwyeDtLVAiX
HxQIuNSohCM8hfFQXOP3NcxnnCoWje5/BWNBRLgbm2oHuO7jFMVVY93J90aiaKUZ
j8dsS7UPwrv9LNqEFhDJ0f28YWRI8WaXUCrV3B/2Ftm+2brKislx2xBbAy/0I+5p
I4koQLRvXYzD/5LZKpaqrpe0XxvzMKLd2L/yLRId1lnHPmw3RjcaznKEp/k1lMxA
VljUb6TWB6yD9i+jHiBGsaMZH7PFWcZ8Mp/P0y1e6ogBhAtS3BfLxAP3SgA2o+ms
MsO/bINzpnIFjzPA31AnvLlT3LDPoULjbp9lIfqut2CMSrkA2N5GNQ/yGSgxOoY0
3RN0bQ4M8tS43hOlZBBp9eZZMAVwKFMvZ+kGd6f3pipFeqVApUJ0KeD7uALdJo5k
dlE0myMHMf2SNihuK9x4gr2Pg8+WiG+XdbQ2YZaZJOy04oanCz5/IqrIR9a0ayOn
k1HZiXJvWvmx0p8es1erGM0An+eiK71fWAn54jZ+mDmFpvBWBSHu91fTyOp0i99f
B/9sBKPQivEKk8hKuc1fILbWmZhPNaJZqbhg5+aBGpFpiSQEg76/QNOJV2dwaQKX
e3XN+Yd5eeFvla+ciYD0XeA3Xn5/6tNitm8xoaMPgBv6hyt7tGj5h2e3RN7u4lC/
09+ozhKEqq1stvifXmc8nkqDG/FQwXAMJ1adt7+dwNanuoFx+tu+kFplcUgv4Y3b
poH3O9hbmexN0j4rbJ9QvWlyq7HjupbGm6ElIl0GYbl/XGv2krhGWidHk7LPRZ9n
6JNprTLPvJVNju1rWZOG7v/r328ffaSYn2bm5jPpQzWX2kCZ0lraTa7Hd9KI8rHN
9LoD6LGIpu83l1Z1CNKTvXiXKkB1Q6HPjzDZyu2Z3lG11jGxr3M+jMRCUBTkvi3n
D5FA+y1FtbUtOsjp9MY/oDsfdt9Q4a9LK+1W/1BJXkrbycwI+E/mMC6wxgKK2izB
aFfk9cOi/oOh+Y5tJdL/FfklTT2hTp8bedNKxpXfv6VG5hNbXkIdu7cS0nNH9yXp
7Ire2dsr5QtojVmB5N0HrsYodzEA6+iZSMYQz3UXkV2d2l1IP/x6NJLXRv30+s2C
FNoZJxmR4yb1ts++O+XLNS9l4ENYzVksPMMQaHfemG4GQTb17Eh9KgKipWqEhjdb
wIytWA34AAqkoDdxGOD5XQQUNNRdY998kzNybBHRA07lDNw/zgD/lvdJpPZ5xx8B
35dyUSO6Sju8l0x6CjcYewdWAGpaKVNSE+IHGyWlApQIYUrgtK/R9tYWDr0Iro91
K8e+aGZahM0h4j3T9ASdGDx4SFD2ubTp38DY7mULyFT5YbL03W3y2gLc2c4EbcTP
aNDNOmLzQNfv0jkuUiLgU/V+2JL+8nurP6Ta2peMX5Zma+f20s25WG2dZJF2EXWx
5d7JEyPkWU4WB1sPmStzCChvSuW5NxU2ijFOE19d6+YYMZ9dp8uVAGcqZcpKIVuh
G78TkhrO0pMXXRFtvDShfvrzu9f8HohdMsO0dMUscr/Zw3mse4P7MCFeaXL5W+l0
qSCeWGrbX5N/rDh91LIMGbbLS6wyQAWL5mGrWKhjRpaZsBc0neHsk12rhDjTLFam
ycefdFXdX/OFchZFTQtL4hB2iKlGcD6vYn0vdIg101DwH/7hjHNJNE9Uoc/u5sP1
he45//aDp4PCT8pKAsdpWVBAlNlqEy7bR36996TqlER9bWmXWYMLaGG+Awj35NY1
NQeUifWRfroEtIUCWqo6Ln4DYYv1D5q6d+iL+HX84HZh7EG9nnfLXSrXkpN9ag8l
cRqgY7TNXZOM0qyN6pMNMUy+FwGDIjmVBzbJAzfVsAZNeHovtzILVxwEtZgFql9E
KE2RfZpjBZDy9nZL3BRqTPO3vaC3flr4lYFouFh6WXEgIOkdyDR1yoAo/FQ2s1Pk
R4yPhfzojw85iWBYHc0RtbFomAwUmsb72VhLWevUwAyXmc8qKuYDEtJNN+1hXciQ
TgL4oVIbyKDRlV43IQ/n/HC+QleXmglMmmecgHfH5r3ygwr1KQUVtJZ2k5qaYqTv
BBO+G5qAUahihKpZbcPQTJlVGF4mgG87CBp2UM34idzbf/nGC63T8+FTnDfKC+qy
vTMTn+SnVAguyKmNPOJUlch27ye7xg6buLE2QEO+Amjf7anTmiwwrVCvGhaqwwUe
fArS0XxJgg3DsoWmq5UJesMCI+BxUpacVEKk7EbvxpZA9pDzMYxOX0VPEAhmiJTw
wZyiDZdnrDTNTJuKgATU1Bn93hxpS23JaW+uXy8kosl5yb+u6YJXKZfLTbrZGBt6
3dSBBrbmy6v6mBSrqpTjJOgRDGNHe/Z6iDfpxyBoaxxQ1jnHVVEzLidBV4isIEY2
nMVR2aKORepw1RBqmVjLNCQdqAWVC3HF2uPNit+BdQNwDyQxuNyUUWg/vv5gp08V
KcaSXpbNNDLFb+lFKU+XbR0k28GjdRWGXQQOJlYbRf4e0toAdIi/Vc4a0IHfgOAf
fJXxBedA68wxN4efOBNrt7UY7G0HRBVtcR5UqNsL8tloiImGIEELNn7HH8wXLcFP
2tR25Ia4od9zhY+a5KiyT9jykA+7rBivLHpn4rSjdABKQZGxNGho5Yp1qhUUYMpP
eLIvbZz2KSrJoxIHq8tV1mswjPL50bhhn2RPiR3jAZnbvJBzrYF6VB71u2B+4qra
iNOa5idVyKu3WBNc6NcLKSFrgbO3m2lcNVGkJgz0GhXspvvoS6z/5A37V+TEKoHh
ql2RFt70gdU1jBJ78+ytb3oHMywmZ4gBE04+nYl/tJEeQ33g1RGCbI9jclWlNa/K
EZiPXN17S2VWtySm1b8ay+jJduPLBt7i86iCUXgvux7cq23mujauQoXWYQAeqH0L
QWJLOFswgRu3G/lkm2iXvyiUPMWPu7qFTDNEUXY5n78PsI6IgT94ygo67WWRC5Fq
cu7b5EGTvL0wiiS7xbRENqQ9rjhXKajhNoeQdpcTrF74zSopgd+DlSN/Z/MuUilx
ncBVhmyvvyzJ8aCkOw6AFY6vX/v8n+e3okWt4tzyZFV+3BJY5AUylqO8yqhj0kOg
Ga8tzaZ3/UJiqAIpPjeKV/dqrlOjYJ4aZVsEnKXyxeQifNhki/lLBSSg2jtj4kZD
1MUSBhK0IMfivLKAYv+l3TiRK6abRGdlM9qTOyL4MTDmz1Pf/IqvmBB7QBFYvyT/
eivbH2AqS9fhQFRZmQs6DjZHCOvBCxbGeCNRNGcTArZQAYVpZvSELGgbTLzMHOIr
sEiO/h11siJFxu8X9o9nllqnI12JeHXthLMmK4wy3yB4sxhealdZXL7Y/ZaNFTCU
U6slsvJaQZ34ja7fKmJGr6sRvvkjmGLHxF0yO/uD4yqu42V8lHob+qM3LyKuAIHz
MnrThoA3nVXdEdjqjvRR3bdpedYMfc7bXwKC/LBzFT0=
`pragma protect end_protected
