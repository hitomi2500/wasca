// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HaAVTSPnYiOjtI7ZmmM2DPuFwJSgk82nMy1tLUlrZuCYgP5IEPQMksUyWvH5OL9F
iTrL8quhCcH7rXdd3V4WAmJRGBIPjtL1CrthfTERHKX8XCEIwSs3UJqH4I8rxTKe
giJSrxM/cEHp+yf2MP0XDmyVFdDfkpLgB3S+/PH+vnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10992)
e41kupcPabPXVd0Tspu7QV6wB8z2evSjr5mfjiY/H7JESXr18cYVgq3s0CUX1TGS
Qbb9daobx67wlKvy9SAKot9MfQyeK959RfCq5/1x49oiRAphxCdJUZLeAAw015DW
c89vo3CNxxMioDsF+VQPFy5hmvYdHrSlgrYITVXFV64XPEYyNirz9Uln9syvVcCn
vWizCp/8yOYdiN+4P/s+J6v+n7/KZn6CS2Gi4gqwKM0XsbwbpYwaWtj5aPmTtLWZ
DyO0iGx/qe97dUcDuQwJRYGI/+d1aVKnZ45McPZ0oboj5/+8yzCQO56JVmLMU7Dv
OnEnQH8tf1kh6rfgmTQf8ojDzFF5EzTU0tJ8GVNc2tBcj57lsdrOJVHsC8uYD93W
vNEX5igSGCdJqiTKlLaHaiurs5aLKFYbRU+BUr59Gqb1LmFy4fLFTPfEt6sZZP3V
eaLphzMUZQ5BQl+u6j0Q8ZkiZHtbFmOpT1ECEs5aheKMy/j0bFmQpXzbgBcgurrg
eC4rgtEVDzc+LtoBadIsbFu5nVKKuxtGAbFoWF6Gc9oG1hDpVhysD2bsqnB3yrQa
ddCpdSWGj61btorHXulmQTv3ayC6D09dPihxrK5JIaX9aLQqw5JhmXrST8lzWEVZ
JeaMlsU4shlLH51uG/y68x3nNjtACHtzBfEb2urjciCvedvzwwqRhBaw3v0Xj9z4
UwJv+g7tzSq/5Jb0TsCZLYfXrrktTLvz3vLhquNwuZSYQ7Y6wQNLb7gROl+Ax2wZ
w3L3Ci4AT/cXAgCXcFECvoZUD5QRWC//PNEMiyNkwU/M914STF/vBUia4rMrjuI5
5jSaCoOJsFTn8YLqi8WzXRL5Zur4ox/U2lV/Eq26sbbrvilqYUIzlAvS7q0HZDXK
1cA6iQjDGQROL60p0SiYroNAIT72r11xuuaBI460IORkqrHJOYMeN0tLEEXWRdGd
2u9KsqxqZAVI1lT6seho+io4PoD5ZmnDwV0ad8oMnSs45kgDZxjFTYWI3ykSvp8i
8el9F6v3UOIzsM+fidxTa5TMtWF9wH8VVHX2uzlytoo+EyWmzQ4tkZn5kqn+l03E
YSCRbynfNARYUNgLtRryAPmadW27Iz7za4cT+2N8XP2XKnSgSUYFJDWoIfntEaXL
dH3E4uXDVPjBeub1HQvwwvgtqInv+LJMDTNTzD7uOnVn4Sp99VqtXzIYu1gKndhQ
ymRBxrkbUaOC8b65KGa7rAdzOw0SNdHLMsDfYha/BgtsvAEw7BoObxx/bjIcbLKH
JWr5XN6GuMUGp7k/NzQ/JBKmNX8BKgF1NlUQME4+MHy8hAwvYxO3gHCLNkRfYfuB
rC6vHzqZ51HbzY7nuMOj5cynEyZC0wQ5YVMDNr4aZuoVZHWRN33AxpmmIrlEtchF
SENRRTuql68OzHwMdaeCsU43clOg6nnZ0nbrcqj2LlN6u8cOxoB5sDicOzAIl0Dm
V2VH6ROLaTODql6K4q/C1yT33JDpk8tXiK4QO70j/T2q8vWL4FYZAU++SSutB5ag
Jev1kYp+Wrgx+nRS/TmqVOg6y9vfeWVUP/hJK7ZJkNP0xtK4DeqluNHflCy2sy0r
D5Ey0CCEJapZFRngREvrnL79pcokNhvp79VWOwpS4emKr2lkRIs1UGHuGe/uEL61
aoNZDrX5p//2pR5YVGiQpIuFXp3SnBcaCPr9ShFsR8yogLBQ/WvvshBfphvjxnQt
+Wi0uEZzB1YKd9NZGRdtdXGrAIXAqZfLzq6PROYBiM2/D1nz3IdHVkdarr1H2EXH
qnG5W7dmE+qj/JfaIY57wnONBj68TBCU1ae/s8gfM1oov7hB2ZYPQOjg37+0hsbV
QedValAUj960KWdwpW4jI57nSEtHqeGj6VnAWBAbgNk7ShXgCE+jxFAABAb2DrMw
irtczFGBBj94z/k3qNHHL2B/9IgacCUK+j2dV4Goj/VRddlLj663taXy2ck0s3p4
Dyv5Ppd3fmkAlZFnu4VtEPEKkAuZ8o3VyqsMILJH0JBiBTeXX8jIPimp5DV4Kbnu
vzd/ECEzco/93kgXmqGuEVzxfdQaqnPc89kAziM8Y0lxc+fj2CIq5Ed9mzqaW3Vf
sPi7pdRAZW7MezAelt24MXNphqj8vuCRK5fDeZCgWIWPAhXTsHDaqxJCiERWLS9G
dwwmF/6o+/jW8YC9OK8VQxO4OMdztO17XAWIXXv5YF58KZC76nHqo1Eln6/uvUfz
aQzn+oX88yxnI/4toaHJn22MUZixqm4HsfqGGca7OKou3SqvneFgC1L6gsmQnQS0
X4MYS0pTmesynodnJZP/ivSLz6p1XJv/kNdRlKRIPtP5gQuymO25o7n+egoU62jJ
AcysfSNtK+qQzatiNUQyRzxJOR0XBS75Sjt1SEPxK8EjIS9R34EeT71+4m8VKnI2
WTYDJ/piry2Y2oKY1ogqzYXvMOnnEVX1boXoE+ThN6eJGlC5XAI0kjWZW1vPYNBM
zOs/Cw0wuMAw+aRvzufjQJRsucmAerXTFH5HoEUOqNIYTrZJzkjQ2ubvWJgE0gkS
x2FSpZ1gSHHoZx+M6NWosxRrrT4qGu+hQuyyTCDu7GdIQtuOBQt+8p6vnyYIZvgV
3nOCqbTVxFZP0ob4X+o+HXFvw8sb+TqdDpsXG0i/zvDQFrr0puZM54p1hisVaoIy
gS9gcwlYqt10vzPT4mOtnyqnHLsBNOtb4CsaFScUDGJgapsjvD2JkXg5X1p5QgtL
JPmuFMIUNuG5kvFE8FLeN6xLmue/AS7ca7kndeCAd8klFj4HhxGHsJ0sxkiMXoHy
PtDEjo7HbF0Lsca+3xqJm0TB5HedXhciQTyZWE+x4YiyTzMYsZB+yaFu4tv4jNxF
JNyee8WuTrhyKo6mni/xDIpCxL4+04wojs65kst9lS1NnbAlc3znZZNElSAx3pdh
+VJDMJHjnCQ/1vWRFcNxUfAlTzsRX2x2vsQZQZ765S3M0gTQ4o+FrJWUPHp4WE3L
Re2JEetxD8KWugZojRbn6COTUFkV1ONNg43UKLwAX1rPIlagFdbrhNR9wk0l6jeT
sBh7mrSoOReOgJ4DkE8nVFegDawQrioTjTKRAvHAA5uFxR6buBXPMt4ksloPSqca
aL+ITIHImYi3fYV02HsVqi8wBKJYM25hS846j0IMmvTRPScVsq+Shl1U/4d7Acqq
+PByC6hvN4JxUcn2sae3QhG3m6F1pVbbD9nHqBWp9eadIFbYiyDlEvTm2AHAtjdZ
bMzqWI0mRE49F4CHG7q0Tizd8dJJ5H6ai+fdtSVylL5u6wdAm1FcYvPmU11l+5hV
+ehRz565GsgNhDxjVsNff0CQScgzj2+gCNVqSTXUz4HdN8+mZqhX1vDqwcSg1ODY
CpJn54SscPM+p04Vfm05BHB9LxcFRgPvJ1IoJUfegM/2Zp2ZWEm/QCzIlqnLwlJC
xVTKBriI3llxNKcKqaZva0ci8O1q495JRYKjvQWgb5fNtVXAmEVBxuXUDwG8vC1R
fzNiwoyzD33rYqy/T3PrEvZEzhlzchSDtO8F/bliMJWmzXCyRHoOvoiFA1OSZB5s
f+R4vlA8ERWmpW6yi/YaMNBHEgGF/gIz9jYfIcyRVAH/F6SK8N45cJHKwUMjLWjE
vf/OG5dCErrk1DztmDll8gJtP69trs7fIMc8Lt0nkinjVhoIP5zVLh6V1TlFwMY8
vt+aD7tCDkTt0/hSGXK32BsD5jIF7SUqvYtJTB0R+L+9cH5EaPZ+FHefbGfGuRqU
+tLlT493vYHX2NNOaMnhqVnFVwJy72NHXsb14qznvR+Rlr2+6nUaJtpj7/5KAx7r
oefm7N4yylj9pU7rLJHNisHr2JFd2bnzrg4+mJooycGK6eZVzP5SOZCjEIRwWDGr
YHkkJyecUpw+oLXf2iRGXeq/wjYI4YJOkuW7YCTzl36h0yX5AIc/66Nk+zp/WOJ/
wpokEZOjVLmgeAS9AKwsWA5vVVCXRB43AdyZGLXC0eKl7l1rklClBnBb/JIb5TnG
lrPETKO9j/kmcmNyeNOCu7VMT+CE65IN0uYK93Cf3C0OQf27xV5aFTVss0xXZkLJ
YhqcrAqmzMOPPALU7IEcUM7Kwd+Iaps06fof2Cs+SLO0YnNUiwklJWNd99EI4Efu
6SyJ6PdVPzEqQtvMuAIgSObK5kg5jRHEgSy8qzP0kj3+ysSU3B132g3010/L4C6z
HAtNAmnaStF6sUkb7he5k0lVpXDcyKfVL8fuYHYeC8lwv4rDaexYPsX2C5MJ8IYt
+sYsRzkMsxqgoTIJeD5poZMD4HaxdbsCJR7ffsOPDW7dyDZF2LjZ7wg2BsOA1rfx
qGYvx9xlT9d0eXIHOC/Te8CEaNKry8+2JwdiW/wtIDOADBSfIShHL3Baod8hHEq1
v/t8TtANG3gZsiK0kniZhh9UpVdazVRtOabP8Cv9cdLB2JQNsEqLkU5S8A+xRzi1
rZqodJFPj0z/xxphKxd/9SWXX3tQbd1iTYyqZbT+q4chPZ+4BpfQk8eZ/r66u/Yo
2wc3MzxqLZFbgXr1bBh1bCZlgTj8hNSv0Zg76d2FcnF3CT8WvCQCYEOLFOofd+K1
+2VWoCJE5zlrMcVHnHspdilM9jP+Q0GH0S/jeDqYctctXPiN48FZpSAp8pm/P+vM
xxLgu41OLkslcxk6S+9kdKadA6gchk1YlHWWepdot2hwwZD1dE8LtwRxF28oe5Qb
z4OjXAsDRhvNaOOhIe460IrJ2rL0b79AwiqtIBIh2Jp9XmtPewDAsFfGOGZ9QF8t
QtANbTyoarEldQUKkqfDbPw1A5FRk7HzXYKEPf2A4ydnV6/XSAnXq65eUNR06lRG
h4V4mA0kC0qiKtVmkTw3shm32v/BPqSWsYs8zm4o/UwAkfJVNkvS6U7Mm1zrJwve
J+lU7zK9JMrfdE+6D1tArHh5JjHNOuO4XtwzTay/jHbq0gE8T/68CrgBxmOH9CyJ
+7agVPP4y15d32TNOxRqOC+rtzbgVWeoUGkc2XLsYf7ykNEFKScViRBS+M2E7WdH
+ytmjW1Xl1gIgJvFMCHqw2Zj8k1Z96y4cmQe5hOp94PrjSyfX+5ADMjxasoXhV0A
OJpdSWeSz8ksHbpRY6RjRtIkbV+KwcvWY1soUmOtpJIluE34hSz1QSz3SSY3NMZE
S27KbvfKky10uu8meJD1fy3jbrQZq9ge/6o7v3dFfLFmwO7vOSTHINxpsWQKeN1U
P2Dwx7pzGsFoWftDLl5+fnkTi398lo4DkNF+I+iMuaX/GhU/pgJTmiXsu3CbyBXQ
ThZrEHTzrQSbXKkfFUzF+cX3cl0Ys5nuf8Yova2hOIauxmG39c5b0hW3qMJAF9nt
hrdzoBe3kWOZy4m6HHdoI6hwdil6bauIBwNwt7KaJtbdrdW6q/s6VL71OtJIFkN5
kUZRgFyJrYsyI23yAC3axiLSbebr/OMdofm6p8WU5ELucG7ybs99HIz+REyuIpAB
IBXUfj/alxDRO5VhH3JM4MBFOMp46qnQiKDRqDTaeAY5f28bMPpX6wBGKV5qoKy3
dVmHBp4C6pQEyZBGpgU/AGuPmxx7fIukCqJ6V7DZ4lx7YKr2EgcbyTX8RCncZz+x
whL24vYZk3llhdsHCBy6empcXX2RjQIhkBmZW/5oInKBwzH81aSWSB/2nUrwyD2Q
w0irJ4EOtrEXMDhiP9Yyr7XVbgg9XPcUlcLZKm6QPSupDqysshjfQ4iCre4AmBm5
hfI1hHf8PZSMW3Etf/7uhjFTQOz11yXqtYRIGLf4/XJ+xOShSwGaPvAX6tEArKQQ
opmjb1xp6/1vlmR6gmZ4QUp6PMfB4jhmV/9zDDVrS4w6hqESY6uisZiaeTLpTGjy
Y20APxdzKh/cNGAAxANlhsSWz/QcRHc78ZXphPqQFFOjO6f8xtXBia8z237vBbbo
5FI3/1ZYxf7H8rVzoodZFo4WMJYRbS8+4Exrk5dF22DDaWi4xqkDN/eYntnH9XcA
OT0ohgu8CNC9JW4U3euouIfd+f8NlmLbVjyWiytArB4xzJY02OGrvaw1qdNzt12F
+BUjrSxgePaYQPweTYyopOSA/6sXcQpSjzpswFOaFhkwVZ0SNdTIdEpXuk+95YiM
vly1KPBAQ3+zSuw5nB1BnilgDRjffinFIdUMxuEsWF65a8ZFNDWoGuBE7/XTBf9W
kxMdmubXL0uh+a9nkXQwzK7F8v4ngWoDlituw9CnSUhJzHAMtTdYvnzamQlvM5Kv
ULNqFgy0wSduofUIex8R70CVfXrpueVHqTPVZCksCxWqzcDGCkiLllTSGwBgdx8s
BjkaxZ3c6IypS61LIZ3O3Vj6QsnuB0wDmrD1XBTxwWGB1F2CbmgW/SXsXPmCfaoU
e+dRDY6YXQgdTyhUaXjr+nOdZ3+Ih164tKqLf8P9gH+cB77i6rS69G/WFb/xJXNs
tS6sgMNJsnUo8bkMKT8BVz0BXf9xDJ91TIsIjJrHdAlrI59vM6stpBdiyOb++9xN
Ir0vJ4IVCmZHFh2+ViVr2AlUVSphQmaPqmfVzrwL2YpDJnC1HmpV+qIeAIwrcK7K
ik5rM7DVOD7CzvdLezQ5ROdsQYqcmCPfDeCEzi22LPHUfUC15IfJiPxIds7M29GW
qCNLPVPZqYdBlKGn0RPnDiVRNAjLfh9IYnkrIMEJb+DB/DyF/5waKYPvrlIv7UVs
07gMlc2NtztmXKkryDMYg+5XiKdzzD7WYrjXDjWbwnKt0AnbRxVc0TndqMiULczK
lXfjIFjXcwzN1SItvOGgMoqt7UJ3+9zqF3FL26uf4c6pBPR0tiAk1ZJw/qTL3O/E
XJnG6/ne5++mRC/LnyUhHioUKHQxiQh2ZK+K5rujudSEoq/KPk8GKmMoePxEpAol
ndl3Vq58pVOWY0x8NUPGlOa+gLJh1aHt42sOCgFyNW/gFq2zNlI7nIhnv5371Upt
wkbsGTG2G7HDy+1ntsPco4l6pW9h+iBsko+uRL5UpN10+j6ZNIJaNx8Rc32LF/ie
pLLg+rZ1tybA4EApRW8rStwF5VJx7O4Ef15zDkAkkCiG/BjDLTQykW2fYdpyNKFb
AqrDY5eczxgL1oB25Oy0OxEzLVK/1aBfgEAyvNyY5UGxqibxG0B0H6irsfhJ7a/o
usQqDi2k9B6Sdm098en3/uKycemIq9NLammy6UlYkho3HIdhMov48eMWhFZqaYtl
TyR7ItscV4iWUxEynUxa5iHTKgojbbBjd+1kEY4DYswuszzE/m1hsAWdGyssiU8Z
kSyyhDqnH+npZ7Jy5YSnIPP3q+wDrKolv1YyMFax3qwGP+3/X0SNQ6YjXEKsazPj
nbUDzHu7hB632oCCuRcn1POwrf0mDtAY7oi8NVTDG3WeJdrA2QHGDF7xwch/xgTK
T2RNw2PUC5g27w+eCHmr4FX8kV9hty0mdY+6+Jl44bAtWFPz9O2RZxHZGsm4eYQy
hf5M6VzWSPDpTUM1G4vI+H/rT3al1WZhQUU1WExXT1n7LAzRW/0RsD+jjMcDs5uJ
z7rr0X9Zqq5jUUYA6JQBKL+xdHFtMz55WHxzX00JoasA42+rrBUu4EMxLGd+IyVH
uCQccz2tpZjHTKQ2vZTvxmD2tDWuN/w8sf8OgRfFXozsbwBOk9zC3Xff0pzAJmlP
XtBM25W9zVPxb1nMnRAmbV0bTKspfNV5gGDxOdPLiN1wOZg85X0u/dKT7EISsaFN
oK6bvDygILAycoBMLur9Fh5/ECWc2+zEUI2IeppvXAtpWhuOHt+UwODGVNjMMQfd
9nwTHB/nYAmPen6Ti+KG0/gCkH0Dpo/iL3HY27JzblFFeLZbe+sEqBEzopY1GpOW
kksW+M3TmaRDI+LfSDruPvspEd5VO/yyw3nW6AGuBOYuU6kmLBopITd+cUKnidMW
UHSN0iH4hvQX/rwHw04OuPVbEHga2gKY7D3zkw2/zwuiE5PmSnzAxJwUvP41oxO1
IZMXQ1Ti9Ogd6B5dVew2imQBBlS3QoOc77Sz5CBkSU7k5Z86m+qKo2SIH9ik+ODJ
q+JwaeuDxVTK7JYl2j++b/BbZ2Si+/tdf5bOmcjogrB4ZKDN5SPsvXjkCnan0A6m
h8doRBPDDqv2lng6MxFaUp2/Rc0KXl2j2WyZZX6kZxayAG7cCHWWflslLXAjF/M/
ejX+muHGJCqzWdWAemN8AYHTMmuhGuarsLpahXNMMff/28zW5cwqkIfKrbbj3acK
hxGURZFlaVAVNdZI0RKgXvQsIzr9yAEXdTueOYOJvcJlQFufRUhpN0AGxmQXMGub
IUXZ3B27v9QmGQRfXfvIYrMllucU9vced+Zbf0JvHXanwVV28NVh4UcGWCSfi6zQ
wfX65KCdMGvt2BdZt0AVTAcF9EeQiwQHbl0L1zLQwvTJbxDlW6GYzcw4VHd4VsTG
ZHrYmEOZytwy/boWwJyJ21uiKc57SL1JDtRR1JJO1f2hVYDioUHM1/JkbN1h47a3
78d0Ava9kkvnpfz0oLkQd3XnGbhh8xAcvJ6bGIply2hBKSjmSkvjEOVS8Dwhmbe+
1/e30FFKix9zLepmLxttBkwIxp8OjIB+m7BbwjOLRfjdZPCSoTz2mIwFVZnrZsQo
VY+g1BbJ10L1Qnifn2n7rBefifIbUB/WFlcYQJkQvk9AAX/qTFKk5Sr3neCzb2ag
po1eaGou/9o5qw/KDmFWNUDgn25wc7G/ZMAqI8J+o8BXWuZVHhIcCRyY4Azaykm8
TqULFLW1/Gu2nMEO1bPyYV0fgzn9OxR1/eyNchkQ3sfOTcQZN4tpRSN7A/UX58Ei
j73rPf6lPTX+oHMS9sb2/pRvfHka5ZGo5SbLXTpwYTQyJo5EIWkILDGBKmRx7rE1
lO6YBx/p71i2pFq/O0v/xmjCQsfcrf6ocKMFCTwJqXrVDOLGBZR8R0CCmOGpFu6c
HNWJsx1QymgTvIHZfB0Y2My6Rf28h6aAaxGAXK4MAGbw1HT1pqknHmZOPXbyJ1QA
M6GrVxUNT3S3/ha0EUipWrdXMKWyP5afeu7pYilYECd0NLAwjj8yh23CvO3GjbX9
JgYYoEEkHvfAD9IM7Dt3BuEY7fOuS397RcGKw/k4xw9BYcMPGOOytJ04SPmpPNtm
kQHSzvIN5kLDYZReY3dZM/QHeCwJ4PMv4WkYF9B2mLC0s3rnYUcGmuP241oMKaW0
7ewcPwPFATv7UGqJ4oDb78aD+FSSm7JXnr2p2n7YTymAKF1sFCadnVvPF2CEkSE9
XvEz8nY80KfC3lMhAXMr6D4fHgJaJEjgcs05VKsLCSnnMH40XWbm8gLz6fb9m0Gb
haB1iiTs6MQqniMDF2OndJ2J0Wg935QFHdVeZwxpAgfwXmiyDLufGLoAGYSk697y
mjTve4fFuoxTQEY/pnmuew6eS6yaNES1l/LGklHGYLPxeePYzcqWcf7of59qPUN2
zx5lvTeA8Z8sfrEvEwdsGO6BZkIdh0P9TwErf+/uqXi2wh9/VXoCXbwUFDId6YH3
0dknhLrJyfYrErP9jCb2nDwwPtwPRMxS0BSkGGinwugXAog9qHlJsK5CKAQGT+Aa
Jp/7JCgP99g9Zlnj3vfW5oSHo3rMFa20JQpNi3HGxNuxoVnHGCHyDOgYSxmDnuuM
P/XjWh0Q8VvqlN9L7TT48Qh908DRLQz+MHbrJMCcml7b6QXOydpwTlplRGcENMl3
ANyu40wJGhcEwc9swT2J8HY14mRHBfDP4BOHtUBuwHny9DGb+Uy3iXWYuUs1aBx5
XBEZFXl5L1aGm/KwIDe3xcL8G/1+XeUAsxVZIpxLQzlNNGvQcHOnIqDzMbR4NCZ+
9zievM+YZIp4W2v/66HB0LhThy71wc2/lMISKSQfHRPwRT38WI4DsP/zHnhMd6H8
1aXrofidF9dQ0Wu0Mi40xIpYELinZtceopLilPOVLHs7RKkixdjjyIfF0dPtS2m3
i8UnkTCQrInEWHcafYVq5z+N7yaHKjxJQJbcV/rrN9+MHR06CLmxKUc4ZHNJ15a6
oc6b1GI/+KMZm+peQ+QkVPgEH83bFlG68YT874TdQvrVxnD4CzkEBZHqA3tcW+VH
pWO+rtbTPOsUwF52mLShp4fnqcvvFwkpWrXUyLRhYnPPUc9wQ1lepkJfUb0k1RGN
g1Elt3Ppow5fbj9HbC/cw22vlzW87jfz+SWfcR+HYDf9zYHKYxj75wV2LH3kTP+l
15rKVSCZRVpKrsdt+lAp0LiVpuRUITX3W9nGw9ydoxf+FFc8pcx6RW0tTlNjs34v
ZFuPlRnNdHIju/uGxYcdsZ+yIod9zA6uoI3JRM+vHpTBD42hkmk7iqMLwERMlPC8
pWyHQXI6aPdSxNelP66OV2hE/JNS1I1iDvuuy8KU67ntDAA9hWfEoVaFOWPboiOh
m6OgA/aX2uuE79CMyy8pUHmvkBhsSGMDzxc/1NRzfYgTDiYv0m5EOenetO6UvCoP
xVOuig4A7n+Kr216F4MH2Tnhi+Vs6xlCwHp8EzytTdqWmX3kYStTGVdE40bTl/KN
UEHItvhjj5uaJvkOWXlNH0pU4fmDDeu5FBvp+CkF3tbW4/0AJ/RosZLHJX8z4sj0
s6VAMaH2cxLjaJaCnlU3lR1JJ2w/CFEA8ThnzrY2GOZX83ivNV8ZK6tpdWx9wXFt
WgVBtpzM8NcGf06Yt2UvOZDdL405MaJ6wAy2ulfkm9Mn8dGRtQU32ruqndBGXva6
KWxNl879zEFFx7JBdTJgRwqLg6hk9bwqaGHKO8j0hWwWUggKLhEA73fQapaRTSFk
pL9G5aYHtgR0qnCE/Jgo2kCd5tWV/Wfv03A6C6BZXrjLLWy/7l5V7uT3qqxnJ0Mz
UjoTtFWMZEqt8yd0nXLMNDrD/a2dJwtOmuw41Xy9rxNIojEP6G6Y/qgl23zRU9/n
sg69SzSG7jaXln7RbqR1/fTBShLcuAzaqzsNLPS/lgKgrnFKVZlqiXl3zFV6fVG5
BscGmOQrXhx6xsct9WgP0KNuzj5yLJOYd+lK5quO7Uvb22v6zSuOnQx5L/nUx9Wz
a5hu43djBgJiIheLF/TFd08K9yrhIJlpYQD83mbJdv3YfkGevgJAkdJK5FQL74pW
dn4AdRNL8xkN1pSGTdHtvM7bEzT2kN+XP9MSQZlcoJ8HaogA+JIOUQmR6MVW98YA
avAO9z+BK+fQNwYFMDetJwOqOdR/aY/ahJf99n1gUAq2gUUIw9UGmSfgN40mF+mS
uEthoTdOK2msWRtpA5xQyfoLFuEi34eVaKBHJLjvV5QVV9zeF4YS8m6uutLM8XNO
Oa8oROGzS19VXdWp5pCl0X5M/an5l/2ot1dut7339cFi707688i0Ek1QeDn9Wz+K
6ZTOdFHBe37MNWS10ZLx0iaQ5nBQIJMSLr3qA/Ymd/f0HN0q7z6RPuWx1yBU3nnF
ToeeoTjT7pkgKFe/dDRk9HtmY+sdGdNH0K/y1GbolTFzKA/XJMpnhyhv07H6O+KK
/BeRyaohZP0RCrgXBRZtfpcfz1nmTB4Zbt4U959Vkc7deOS2yhMQPrZ24aY6Hzjs
KeBPvouXVvYiPrBi+P3qfMWIPbKzBBR8Pplfg690hyHgiiAg0iq3E+7GO8qo8LhH
2XcRVkG69so7q3Wi/yFE82WSiqKyhi7x5X0lgD85VbFkHl00FUPOi45NxywDqApu
YAdXKDmk79VgqGOX7+nAviyfsm035nDX3x3oCtef3A+OGM217bsRzXjACMS4RwgZ
TDyj/GbKT/vHWmcEDDV1oca6oVIGx1KdrNljIslJzcemn+CBr/A8pR1v+lwTJ0KZ
wCTYVVlynidWtP4/mL335QIDJ+6v6huG827E/oPs6PfsHboOwZ20WN8D2gg0G6mu
yFg3g9Wc3y5xhKKoo7TRl9pWdPqLGct58+eV4y8JajN9jH9d02SmOc3lNyX7k9LT
HD9VmKI5cGPLAcC3UW8NsEOkDvc3SKb5r2N3i0wFuPbDukN4kej0Ir+M+gUU948J
Hblx8ejbbyppYvg75JMJatXySBbme4UklzCJSzafftddWDwq/PgE9auVUYe1D/Je
7cCgqE3TJ/F7KNYqNWUwyzed8rAC02lSs93bVysUiu/XkFfLMlQ6cklZO5mkVd9I
64atnVCV0zUMIcugs8jyHjiVCz9Lzz1XLxFV+LZCEsKbxXCLygYj1DQChmkyqGTM
RjMB5weWAxi52qYtQ9LigQ0MF6qd21mRCWG0NiBxlnWUZaKYA3X8kiqiBNbUYLGE
yIMaEN00Q+aR33nAjtRksitjPFvIsIQPLJ+2CKp1EYdYBM6ARlhWqwq5f/GHVbVq
vaxxZU/YBLshn+bYAP65SwuBSa48fMeKfKa33HKurhnS0AnW985dSZnByw3PVmpV
AkDcOfap+7QoETup2fscWP1JiuAIYHxg4CVtyuBNJRjeRwPI6RXE/E/mTnPaIfsr
/2tlEZVo44lANXKJBh355Yhc67kGk7FOWSAPucq3rvea7u+gORgpdeljO58CI1Wt
n5Xrhq/4KhmTzLReWs8x9VaRt1wAIt3ra3whWoGAsomgHCe9tLlU+7APKRbJt6NB
iBNmwt2VBq3gqjCn538HlXSVsWOQeO4EiRBNbiKdJoXKQBB/EpBz8zqi/SSc4tll
a+sC1IukyPhvfq0Mqme37HddBH6XAFOvDAo/IbW2iyY6DgM/g4Xz5qtotoyVbqRR
78z5EK+dOSWZWPaOctGqVjHkgIUR+B1MK8Pd/Vc8Tjbe2/u3Du62yUc20/9maluQ
AvKLQYsIP07t/pGRRlokaOhoIjXxLHiWohZFGSdLaCI8fBnUN0vhoTKwjjiPxMHI
dsHh2R7QObB3g9WzxzYy+BqDFR/JFY4n6S2oobkVClj7YfjagyvQI2NaotqXF1G6
fn+8IkJoYOxE7/iCOxBDf0WbRQmcAHOcpoy1hn+Qz6KV+eNG3QGPoUPs9Xsqehn5
UXuagDNND4y4FuHArUB4c0VgWRC8khj92Mv8Fw9Aj2TfVeWKcPl8lZw/OltDkKNj
kpe3ofiT2KzJcKA7/uWjFgJNjb8Zzyd381GRfCxIxHoi1b/wsrmlPBZMsrlZHAuP
9AWjiGOm5nGghhVyrUxw7n5sMA/SCOlm4bPkd4swkZiwgue7ByVe+fmehtySeyfe
81e+b3mjCCozvu5EmbuJQenxmWzzO+17V+WsfdjUa9I0w6y4vDajDvTl0gahMkwL
vvyeI9Jh72isyFuGw+ncArqsu1vZ5nvr62HFZKU8fa9tOPyvV/xrReZuiZ6c+qg2
5vSQC89jWEzJOyJduAKIpaFJJmtvL3XR2uGT/c0I9JTKIH5BBoyLFsyrdmK49Nva
X+LlkImtrg6WR/Cz8/vbzmH1PeV496+87EyZJ3ZDbeWWr7RNuBWtI2fHm4brgrKI
zhc32GfdtTlN9aZZFxE775fbPk3hmB/vUPRtjoT+TzIS1/3qrrvIuHgIWp8XcGkl
Nk/64EAR67Rqpa91kttSz9DgVnCBkrb05B4gCsz77LTK8s1ZjwFsJO1iLw6pUkii
utazlO74QxhYWOjNk5H/3o2U/igUWYHLVtn2Gg4pXjOiBZ4O9VvmHDZTNCl8A0m2
ydqUZK2GEW7ptWDJ59LVJ1etDb1pFK0r1HwGMvTGA4RF2olHucGzTBebSTPNuowq
LF7gVT6F8nIhQCf45H909oytmWnJGAvaBJguAqHV4PhCOdMjCBlJnX6ot/+8GDxj
7NwuqnFTvEDjOIYhJT98aod4GNoAHXVHs7hVlOyK0eIVH20DSkREdrG8G0fXMCHn
VkQnPVUUpSRXrSzrDDTNJouyjVkBWp2ZB2hPRdZG7SHVilEhmtVVcBhhSYJQLQS4
0EdM5+m8FLZtdHMdjuRP7IKp56uNxVEwRa4r/9R/u01uay23ZhLkMmYWNx8hjqBH
HQiydf6LUE49pOHMnaq5/Bb5XBtus3XJ4r7ynUyrRZWMmslj0Ybu+wbBmruwyJnZ
P26QPkCISTHb47WPuV1j77JzlWflz75F79end2pNq7ju+yQA2shLQROp34BHc3fF
1tSIdts/SNoRqprztnNwtCTED8Gv4nr6yacha2EdZ2pcZ+kXSAu/45oTgpwF74WP
4kBbVOkZ683+K21fK5NxxTiNb9B5WRLHDRNooV7UanutMri9BLx+A7HeqDxSS7ke
BReOXtmvPEzaggO8Jasj88BJUFg0vYUOLkhq4Ee6NAisAMIIflh+o6ZIW2ykn2Re
yIxlW+VA7LKg+hDny004rjTqfLgEt9b/TKrXMCgJ3yXoWJGRkTNzHDXp69PH7frO
MhcyczhlkP8/qTgUZ43cohNtvt8fa6F0bW9HciC3+r2vSCy9r4M4VOxAoHhjuSdl
E5xuM8li/kJzUVC7AbJO2c2xXdjLC+W3y3aZnGmDMle1D9S6BaHh4Z/CtDwXJtJZ
r8TZJDruRh7OjE8dKs1fU+zrVCjmzRXnE5zrNuTLjlGWP88GbUHDaNRUueV2fV6w
Yverz1FvtnnZwFr3i9+mXZ0tBXGw8LOji6G+oBnXQ9gjX4H+1CJD9g3g9W3mk/Lm
gINGg2S5hRe0zdf9hysexpC+wFdv9WoXoKjym7avwivT0cdkljabtGizQplp2SVv
`pragma protect end_protected
