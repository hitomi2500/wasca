// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bTiCLdR1POe2qE62GURfjBMRMXKr4aO5PHR/cM0yQX1/efx7yJQN+86/AVjTi+MouNsJwe5TDgqz
J4Ay7XdDhmmOkToBapyP6MUOKTeYJFRVioovjmZ4vt7BnzWDBz5q0b3d8u+HdWca7w8bC/kZxxKD
NHcVvUHUKuC3Z0l08EojEaozVpgp+ck/4rjuhUGo3AaveE9QOd/B9mvlZKtwBMn6t5U6rp8I8HjM
Hpmkf1W8hb/0uhjblgrvQd8R8+9zUpYEHn28jtyDT1p45I7gHzz9gFqdW4XOWqoT5gwNRvmDodQD
W5kyJi7RBZ7eOxSpqzi6mfpU/RB7DdSdlDqD8g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
2TcPRLpMRIUDRCrQ+hTlyuvmXKUdYOMlCk3rdMRFHD9qzlfRlBULM4sFnBtkLKKDUzXDRPSHhlxk
veABc0BaJtAvsWyRTac/4mVuJXvXLxLrX7OE5uANjmwFvJXNz5ywJMuf/DsMzV121a/8wWgcXfkX
3oHJ5lh+aDYcFiAEh518WtrMnvU4/A7B9Qo7txSbQ3PWedCwyQ3kXad+/MJUlH6JwoNiJVnCk2If
IHwogPu/NMrCjXthh2M8zKYywp77l91ajiwDWqVtP8ajw88DLIhtDpeurRClaM0qEuNOtQpVDRB4
nXvw9hco6onGpH9hYVkUETzR3HHiAdVRdSr9iAu10unBWSTVxIWrbeMrLrmWgyaq39jYw4LC4/pg
56eGOnnygs1MzaCLJWit4MyUFCqbS3VHj6x2jYCOAwLpwMWqnhiPZ+Jc1N699MOQSkZP6QVelREQ
9wPiyCJE2tC8WnEgoBYcweUxpW0ulDrmVB7h6LnAvJEVv+jJhJT0lcTJ+fIliAr95nW95DMUGf8d
UrzIFVaWb84S3uTDXivAxw7nts0RYVpUjCqFe73m7jBHtP8pZPjzX/dykGwkr/ky6QwpPBwhdsUF
4KmSEFHb0/IY3H7fntLajvspr9bwLExNyQ7hhXSXJhB9G25JjoZqPO5F5JcP7ghq/t7rFUIXXWXK
WXHAzXpUNUNKsZn0e772TDlx+43xSfqLA1N6Zsjj475LhJ6yWO5FyAwcVBCarRDfdGbN3mQnomNw
tRYkCoQXhUQ7fuGvHhZWw9YcbrIc/IIxf7eBaNS9Bsj+X5hNrBcbbjWJQ+GcZc62upVnkbIDR53h
YngKyVXpmgcJqRJUBuZ+Dls340AgYnRkvwnLFBkO5iJM/CoH4t2+lbolWs+thxl7QxV20R+INDuK
z23c7QtmoHunBsX3UwDV6XIkqY6gqSjtz1NOE4mo2PG/qXdt06OgdZ1gFwk++WjV4Z2z7OcpCfV+
qZsLkttNtsk4OQJ56NcgZarJPRuElZHtgnqfeav76Ml1hNQJS86+s28Ej8vYUS7/Kuvl0AZu1hyG
KUKDNgYlYkMCTUexR9YW5sjWGWTpRYxcvANSzeOuWV2K2p9KYD+8D2HLvMEalTuA7e7XBcJun/Nl
/iZlDvbyirFsZx2prk1/6dz1aqZ2fpCxKwhLR+ZL8I0qJzSrswmKmdB08StNQujjwRx0qLROv234
8gWAVkJNqAPSZNFSEGUPmGURZYlRHZYFkG5uv0a+/l7aXMcOLwVBDvA46MjKp0XcSxIxrrxGY/w+
zNWKCsr/xf+R2Nv4IiHPSLwf/LIsAjAMT74UD9euCu06ZrKgGNswTIBRx+Q5Ww0VrEKSILav6j6Q
ugEiL19HOOUvCx0UphX6D21vXNXkYjDXhk4KSuHhXEs9j+k40DlQF/cWx+xf1vsG/D3EuqdS2PSG
usXCcAM1vT8uvmubhJ5Ipj8Vynt8Up7mXu+mR4thR3OPqakPCA70q1tpbp/L3rDeyrYSu8rVRaqD
F3F6u4llVJHyoE7v+N2/+9h7L5+bW3CoC6bKgUZYiDrHctvblL4JnXKeHWy9R682JycWV+tGu0ID
85qvl0T358T5epdoA7RsRjJUm3HtwZpHFsqmeegGQPIVERe1+AEdlDW2xeyiVmGQBmFARB4UsVMW
RB9aIuqwzDBQbaeqx+wZAyVAsOf63MmYAygKMiNbmTmCFEhwEccg0nr/L8pqrwgAKutgA5RUPhw1
GA9EEsZMXQoYk6E3MRZNZJOG4N0wgPy6s8s48dDGpCJTiLgKiqpWhqmrLu2UkH79oOJd3YvgeAah
GvJwXXE4N0J7yQ+NQPqrnKUUrYeWSA89l1JV1E72opJDgM9Pqtfv/7j9zspIgmTDy92gTBPr7Q/9
jnRNs28v9CzGPPOX00oeI16br0HJYi0h8xW1I9SjUFqObUa/vrCEs2DYV1B8iTghFMoy+/1sb9ei
oo+1MmPlIgy8pB+/HPwnuLWndUR07hGdysinXsCzsAfFLC0B8ZNVnQFElHAU81rPS1G4ZdM4Sl7r
rNRi+ZapsuUS0maQecms1t4/FK066BkAK5m6IumgNObXTDpxrJXHYGtFRGcvC0GRpSaDMspXkwEk
EyagVDZdZY8jzDT7/kQO7gz0IZRsseozBDd16ZRC9tR7AQwp/sMyLskRZGeuCbe1Fe7dlbNXZwF2
465/fWUzEfx2m2g3Zr+Rq7Vho/5jNAPz6Q28Uso8/WrV9e/5aBXv0l2/1A+A+owAqD3dyNvCH2Ig
G8cZ8mq/farB6uorYm5fNW+c/iLH3LZNnw1QSxL0AJtYdshS/6B8iCaZYsxPQvC8e0wuYvFY0ymt
8KjRjwcsSTwnJBuo81U4/6Ds00PuMTWZpchln8v11YXPASt3coIvNq7hs3VRAov3TIWQiTZyGQx9
FRi8Y3J2fvfiw/Wlr6Xp1zp0ln9/Xv95Vx++1hwsOgR3xMaAsWBUevrOujPMcO1QFy+5OxxpZzN/
gGzXZC0IjrRllyFdvSleNZiGQNv1RphfB0yQo3xSBelRn7o9+ezGu/ypD1FVPzOhXH3jZjx+ZRUP
szyOVW6ErZqgZnehDKUD4Ry3QlDiq/lek6XjaKhu/dTfuBku9zod5RuMBwqFrKGYbcxHNwdosk1j
FAIMadVaOBPevTq4p2UKn7YgvTEUFOfYrAlnK6zi4LNVOiQEGPzSmbB5p82JOdH/5bijQLkEB5YC
rVF4SMMJoa/Zsrhg+g6zCzwptwhGQ7C4XWa862kfBb1kMcqXTE3Na+pWjMRppDNYGHUnYDrUfv1/
ddww0DhmTlhHuiToD3I44FBfJGWRq7Eh0CdRR5JjNZh22kk5PQpNDxlylsBSL4NeGQWOfcwmUQ3O
6op+Umfp92Doq9qIOanaBCzuaMRc34aplo7m7tsUgb3QPm7xi4UYka4QYhjv3DDu51NYas86PpwV
Q1PlpQ/mwuHhHEx8Fr2vNd9CY4DmelD0KkVcorV9pUJyK8sxe81c/ABzeN5+jJg8Ez+R+DeOCyda
YEDtUEPXyMKNdi8HU5jX+uEbqqP6XE5bQOy4o8N9MGTZadbcjanrHmh8rvuhPhk4KL5HUC6scTXe
J3/QNDF8kkEMAj4ZCzO6PeD5jiSfM/f7ypAfW9+Zz6WnycXYWcPY8PdEEI/hjtMJiAb6p+JQ9YGS
GyZSwzjzI83VBM3TIB4DxAmv8tgK1qrOTVi2tAxwH8dUn2l4M0TISBim/4/0OPbbQpnOpcuU2fi/
1KsrG6LpNXwC6udAkHPQHgp3zQnhbYN9lr+E+2RlUEPPWEMegA0Ej2r93Z9hYDwip46DGAiFmZmF
1pqC1x1/xkPXj5N9N9UbNKz2FcxGHQg0ZKgFpcqpkDGEj3Km+ADmkpcbrklDuFTlzvbpTkysWvxU
ykwU9mzuiFP+wsdW3HDY3Q4yAO3UTuQW3JVbEnnFfGA+oX6BqTkDWGcvWEA5956yBeOfQZD4pxH4
YG7LdTF2EcU1m7uFVi7sO4gg2tIQO0UfZ+X4bJommTwMi++otJ0g2lVbkAPXPNrHwO+4TnPW8gIH
F6ARY03xKX4uwUZyRb+v7MENNCQXzTcUjvAAFBo1fgo7BDT8c0MtFucIpTqvpgVu4B4ns39HDCtY
GvQEUsgs3C9yLOFtuMd9Zz0R7rDBVHDUKGY6FIfcJ0fbLGxmMCyEqRH6/d7x4/fs1mqDwcofPSqC
di0OZQSjY5UxzVhzamX02G/QcHMgQ0RZF2cQZLGIwdBLoX/FmdM8ColH18HwfupeR100FaeL3ha3
ldRh3pomqQ+oinBcqDRYZbskye5SKxfLy/J/S1f5HGwB4cP74RBqLj8WTUvOv9IxOmJUtiA14pmy
RL/sbO6jIcoQ4ESCVyrLtTOHGNWnGdipRrf7io7rqvldNkHHcfLI5MjzX4Dthf50l3cI5CmpdS8n
ntIQadC5yd/hsZTvbaJAJxO2JFyvHPnNlPSIvj6DSItXRXYPfrrVSGwH0Qy+ej9FTaQpSjoUIrkw
AWOCiWf0yUCdaLsr0284J6t1eody618vJA7VA3XZuIIbsqukXlHP+5vrnkmv7miCC+ucuf12QKsC
EvkSajsb5ANu/D6WJfg4YMpr1yKY9CDsBYj9zecLJTNAJjeqE5Yqn2UCB17f4rio1ybrzY1LP5KF
JCHhbsU4Xv38WD8LoJz+alW+pPQPrnfD/U4zEhmyJb45WF24uj0+4jtJwZpvXk657DVXImKrGZiw
pb2WYbKdlsWzMf3bYffAzWQhFPMefXw2b5cZG93l+Y9aeiXPTGQVRDvvWXTspcQsdMUctVXxdtZR
MLcHvU4vE/G6EF2w/0jcRaMuaUb7vbEgkR+jL1tAp5TUvPFdXxIpvaFDztHNgfbuODqlDWWm3XUn
c7He06cteolIlM3VsYDkbuIDBiMtPccvvQ0+KA+nXrJ/rilFfllN2FkQSvukS+zzI9CW1I6ERnzG
hBCs+akRUhE6uAFZ94SzXoVcXXr+c1oZPRB5Gsh47/UM34B8l6hqTQK9yRNIT3mB+mvM8YPnIiqT
3FYQZllgKvZPzr64KWomDwbZ5ouYeahVXYdVAS2N+8M4oIGiphkZJJ3eC9tEbW/fqB4GdNAZ3i8s
CcaFQcQ79lz74sdUoAvfqXBmFbC6XAGxETvu0UilIovISvNbKY6EkFuQI51UJ5QHV8sqEdt3Nwcw
JHI1WVnmZtEhcIjhdAKzYOFLDjf/7DabCHtwiNdHlQklfvJajdx2Kv2/R/5bf0z6OdhU4ntjHNaT
KER16eU/3Adm8V1prCij5zz49B4t2hsnRPsBpY4l3eISnElG3ba0Klm5EDcpDICmNhobNrWMcTpp
CaB3dU1t/vEFB8qt/Gx77DsXSCFPjZQP/uWPZs7vYkBBWpCc4O2gy4GeF1MWGZFbMEEXkrMFBLEX
Sa4NaZIRhwuR/6w2o2FvAEZiFUuGiL1ZaBd6b9c+/tOefvRz0UbqMD9WRpG3Xhj47FsTWO6In9uk
7nQZ1zclqG9F8XyrR7nmhSXKf/i9n1PfI4IpEDif3UqLnJhyGpM86QBUHcIiGrBcQtugbPk+o8fc
4olOrRrC/wZVH92vL7xPfHQTJJERLBH1CDRYMbeh3jZT6y3sC3uizdmyGlEhnahzVqZgGm8yqAK3
k0xryz/8yjp1izscuwP62PQGP0mcxZ1JUJx0FyT0S8w7FtOzFFqn7zS5CK/WqEP+m3Vw0+6cZsc+
QGROnhBfuf840G90euee0QtZ/qQar1ieL4zVABcpT6uMfJjz3C+iQN/XA/RuYjjRdpXbaJos5J0a
Pigu3ciL85b/7tJV2wofAPIxaaCNSgCKFioAZiyoZm19NxXCVJ5HP1M0azZ1VHmT+m85ywGBt+Ir
QMdnY8hpUk13/AQFRZ4SXTDJjiaUHmAQ4ZQM5BSahw+GLROQZUeSx1kGom/WNHKtJ31AP69dIxqm
Cj09Y0zFWBKMdgU8c1C//I1O7lgAVg6sI7qE3QofdRTl1F1b5H0k7M9Cs+qsUxyImAGR+cuXTkIE
V7kRe7QvaGrOQFbZTfwWn9VWvrF69dX3LH7IBUzODbs0kembRHalTwIs7g9URxX+/URJ//CY9x8+
xr5o+112izv7AGJNdKH8KxTtxaRhrUGwZoOW+52hXy2lkD1zIYStHtD/821sIUW0T0pEe6v2zM+G
5AdLeulVJ7T8ky9DSsnjjPqLD8i3n6LzWoK6ISsvIvlYSzclftB7CVRzJFC6dVMeEgZu/dgMGRX7
MFppRax+A1IVsjyrAqAW05pzYXmtpxxZUKXulymX4hXGhZ8RNNoWCfY4Xrm2XC7bgMDBSftJRJsd
7MwxoqXKtv9eeQMclaNvwGTsY+lT/APC0e6iIu9s5q75+zfOsN6ojxod+EFEtD6FIk2cYDUgNYX7
9qxL6dHY6T9R7TFTDkydDVzfvxdJSFejWsSvNhSqz/pwv45Ujj+AlGOFRCAOTwP9xtHqVFXx8bsA
eeR7S8XuVbi//ektMbfbHvMaEMHuZFNbkv9yNng3hyn0wZ5Mo1oEh7JazcG9IVnarHO9qgU+krBJ
frw6n8naj5cGFrD0DhnCCsvscLnLBR3OsTvBjktIlrMz0ic6l0lbmS3MVlBYQ6F8YBSlXKFPvAKu
hEsRVsOPp6lbZqON+AuzjW5ZjbWfozwrnHyXtVnfBFBLtPhrlMGF0P690fk4H/15nfkz3MDkr18V
p/oVvTH6KeV5sNQk5+i9uIdzoZTwm1wIQeaOCl/PD2Jnjpf04mRzwjzwD7ZLzowUGn7kk5w2gwlA
clJcYUwKWJI6gGBlWD6zsx9ynfeLB8a5YXNR2J1exlkBT5XTZPRMfyjFyf2Fd1ufgQwlKqkOLVOM
QQ7FywnZ9l6/eqowl9A2/iQW1XS6yg4bGexagmiE11kId0ao3/mxrFS/mPbqglOwKmaE7t8IiK1u
J830nQFydONz9o4LgC9RcKIXoLq5VBRE99h29+1lLl3pFrdOxZIL0QXcV2zc+AofZgoqWDbIrX6/
/YnjH+rZl6hM30C1DdE8mMsdNQ134r236KalI/eYhYusNlsDf2e8+yzl2S8WR4rAsElmf5pseXiy
XCrLwETDwYHOwCElDcZ/EjKixrt0rWJmBD6QNJxVxmOExBG84uSWUF3KCA5yf3XEexublHG/SmZn
Xxj9RzGNY+ZnYcPy8E2Q/CKvok7F/fUTTaHwrdjUw2uwzkpnw7OyQlTlN/lyTIJc+5SOECp8iiBI
qH/c28U3nL6uR+WBsJKatP7KX/JSADw7GxEIrnWdBzCKh0/ME7G1/VIIM8c5zAr01azNjN6l4f/g
OcCC5ZY0BIvW92vUvEPW9+e242fl1r8laSn2pHzToeJpNo7m14n26iez0v6V05WbdOPA2nG8TKFz
Mr6KGiFWCD7cpU5ANVinGybjGjQSMMa2Dqg6kLQH6RSuAcXRqWhSsUZe1B06igvxhki7DdWFCbgI
+sdiAAhrpW5odixig19k1zM8bVvlC6ZX/5dgD69TrsAt+WyHTs5xpOkk0aXhLRzjSKe7PaAZT6xd
N/sZ4qFptlWGYKNvsXWcM5F4tIh5qoGw7T0hO+qinh44ysnSAW3PbHtNVBAGGHOOgR/nl96bGmgA
0TNYR/H811Bojzo9J9/4/8pXtUqw3gvqSg7u0k1O7k6tNuXAonNJP4AeoVR6yOQnkS7sL/BTL11D
OYm7HdBP8taImeZ8g9aoR+O1p5c/AlzEJhd/DBMA4JiJzg39tI8eGmZPRFpu+pR1vEqv4Uol+hTm
+3gO2nh0yZkVBLrmF+UHbLoarx34lEViPVgrq/qilRA8o4RvrLOPUhFAsJiVwENIPuPcrnaZPVsA
Fgpm7Z2JPJEgIq8+tG9FZLTPiIlCgJN7unwG3a2GCYiP3sxcfeWEK3nD4ahSAJMWdbjQkMvw90x7
2eg2xucCo9o5pm7H715oDYEGauH8OwHaE081/km3zEIsXvhxwNkucB3ggLz5yxkf3X5LEUXOBs8y
Wk3Er7dc66fNgo3TPlb7EWN3tEjIljSdDhT8YFLW3wN4Yg15IKwoZ71Ai6nl+ZuwcAIBsXapWEjK
oceQ5BFRY2UmRuwL6cBSpFsTR0Z0mIIBBSLZqwsAVypdyiZ2ze1U9hTQIko6R6phjDCT0fDTjcSA
HR+Z+2OYJH30o65JjckrbeUfaCEKkIMU6WfxwEbiNaoW//UwtJattAB1voY8fwTCniepduuYyEr8
GfM++IUUF8bp17l/8Hanw9CXwGUUfc456CG0snoY+1/Bsp85xTCSZbA/11RGDuXq/4ky0hjdkDoM
RIUeZql/VXzS/BdyQuewhZPnUjhJJEUjDXBD9VhtxzdE1tyuHPqPFJg18MMwVp0vHirNLhhKx+Lf
FGumS1fsd0OBtUWFYIWEaYc/FNSEmHJXSzZMYni3k+YEzwLNO2agjeOIaFI4ZMBtepikUIzv5hCl
sDq5C31IN6bsJCXfcepFjiVu9Kv7vB31hY014fT+mksHpUlAIu3IWfk5DROtOpOsM0d6nj3R+Tgd
HdoP3KPur9zvUBoUCqnFS3f+PEBmvZfzPz51oviKAdc9lpZR/Dt0SMLwMfk2o+RqL+a9hUUrjTDV
Z3qInCS+DA/HD11+BRRymRSKWu0lpKkuC/9yZjeW17oDMqhiH8G3E0X5E7Aacvuz2m4rsNC38Nw3
VXMvDIh8d6rCGtJKFNsRTnICxmzhq0tcjpoL+mRk2Y916xkg+5yS3rg36ODo0RFLorlRgry4p+qT
7kUNkt1aYVrR/QwlJZZvWLZXslyiiB/x/TN2p1T/QUr9KyTxBIt8oHobkcE7nU+34cO1IBIxfiI8
WSI9peQQjYayz4k2NmQIKZ7OTQMGobCCvl6TiyFj8GbPspGGo5NDiRLJehD+4jlsWRu0/58WBgxj
LJpjZ22OooCovJORxIG2STUyN0GmEbpWehgqhzDRTKjegwbteQTzwIhwGPI6PAZFruJDwQmP8XtL
ynuRR6+/f6GLAucYeYahT0qVBkaM6cKrTPRRSZ6xAVHfK/VGOeD4JTLwkdt82Gubi9hxQZHGkEI/
JfMPOieKFfXp0E5tbcDBWe1AlVTRoRIM4V7NwAjiEZukC0bibPobHZ/eyNIYZ1eHrNS+ToL79CaN
+MaCx+u6wdOBSmf1A2c5l5Bp80bC9Lty7YTUXpGQ5wGDfaL0n9LPCQk6PKUlqkIslq7Nc1RJOVz4
UN07Gs1E/K811yHClcJylfQGsjbn+g0c3KG5QKr3Yuf2wuZm903o0lviV8YniUWOJ7y930sb7b95
OWkOc7SiT4eeY7qnwdk9m0wlUgktbA2GgOH5DthHZdJNMRu3RsaHR6puaebap9w5SQAJA/1AyJga
9JYngJrrW+XWG13pL37EwYBEBsDbvmJlzHUrMhBVWlTo/3Ka1+cCLMx+fadyYp0e80jd2wu0kY2M
ElJr0pfBmwdRiEpCICgaNkWXggE2noGbJdUIl5hi8vzj0EuHwHerOq/EO1o0TEeNyY6Hsju/ZoLo
Xp+CERrXrISqqyEUKVqsIoUiQZf6bBdyF9uCtdymKrLdsUKlbICIejw/8hgbJ3irTDpUkE17qr1F
34AAWG8KMobC/ozH4RtYpq3GRtU9ylkzMqDoGuazImlYba0Xpew+63cuhfdEh5uUYI/slv5cqTMd
8Q9MwHEXWxEJJSAHnyfC3e6T/RJCzcrRgykmjyuyvL1E5GZE3xHgjBntaR0QgyrchtZKImqUVkCG
CPBo/cOemTV2JAMLYSjo3fRLhCvcSzzbTUnxc6QttNjEt8mX5fJepkLDJPZ3lulEOF5UZqzuQzK1
aQZSN+Zu/wufySOn5GnB47zAxvUm4cl9byleJq2ZG4m1Buk4I3ENnny3x8Z6yuz/Q9MGBEi2yMj+
XzY3ACLA75oT1f+UINYtNh7ai0v7XeTmvsCXq2ncbrbFsNPt8RjTWyMXUCzv4ohNeW7ZtR+Q5pXr
7MUCX+2aNVEMt/yo06ejVElEmLtY9sN2h1zC7EheFizGZ/QqJGlTfx63a60DPW6OoBaBphrxGHle
TfROgGm+58pE3y4bAEOOnJkNTCJbBNFw6/f8ORJ7NFydlqyjCp4E58VKYWpcGK63Xf/5GonGpsY+
5rfv2Y3agXyIcSIyUnTwgXNWGUmQnkICn3E9JWOa3c/93RoZV3UJgEiFVOc98NgXSiuYob4ma2t8
njddUvDKRtuGBhkgIFgzNjk/APdn+SweN9z9SsjJvwkTtP3sII+H8yfbOBRi+PG6rg/GyWvBBt8i
0+O3tdl/j3vqCR1Z028n6APQ7r0A3wfeTf3PdzTgeHf1wMjWI4kJP2A+8SmOAELe9wUkNp5PDMOT
u6NDIwuW6aFkaBSzy1ri7I6FAy4QNImk+MDpe2Qv9+VlVQyFyANeLXCOj4dggzVQNudElcJphxtE
oTBrhPYfiq3Gkk8BdjrBve/SY+VLR6FBYADusAd5NCQITqj7HBDTN8mqlFTkiOLoi1zv0QoSmtiY
7jrtxSgyCX+rWZ0NNTYAUGQ2BH4yLcU9fBKz0qmt+NtQ/ZA75rRg/b2LcQad2iYwJFPO4Lj3RB+r
QsC8f6hHQy2k8G+RDiTvBobrlHSCYQyu+c3QIRmFGeRBY04ql0Gnd7ohyOwu1SxJPCWdFJXO++5u
0f4ZKIsWMbh+cth4Qdjknnt2ytCAMhZZwZ7rwh8drPYksdNe07cRwEDykuFwXSO8e/ImCTQV0k6H
OxPIaCmefZSGgrhVI+Tvc/QZxS4UQgYs2LcX1F0W/kKhIq0tMp/6YvfajgCr8U2tGifADhQc9Yvj
2JK37XwPR+RR5CE+WTttIamVkEJAj6Fw0Uyj0II1ZgtxNZt36CVmwWFl/IFR2sB+g/sLuSWHNsRi
RREQ/zBipNm21PbsBgoNZ57CQ3xwfU1YhtnzRmI2xPvL48QYrDLK2SNS+8/Ny72qBO8qo41UUO5s
3HSoMTLL/hd+i8S8x2v4QDuGOYoDqUdMqkADLL5dzLOEGPuKPT3KKxvow0I5m3A428tAxFq1/r1l
5s75sqIrcc6gW9BzUaLP6p1qzRlJJ2bYZWuqBVt9n/UOknJADB9TFODKfuaKPPm6HUOkfhlUvHRm
HIBFqH7EV+QqR3zIMH5mRZh7Xi3X9MO1nqlT0g2JbKGPzJDcUieqNTZHmtJ7UDmp0toQSZZW2ly7
pBcj3WMqaU73/5+L3v7k5wmueXKH0ob+EHvcRhMxQGCWsy5zd3n0GdNpYe8LUeprRszTXinjzJ/h
jpuuTJF4IDZxvweIL/f0RfOW5saPHDXEIWkxkt3eDrsOJ7kZq0SnAWY8/nEHcLGx08vPOdSZct9I
SGcBm652xltRQYWrFKFTVzRcP6W/15heOVfTRpI1Nt685PeArFIZ6DEhyEJXljrYNeo6qTp75XYy
OaJo+Z/30Y1LSJWQiGJHTf7673jrmA2G6pvsGgPUWCDHMRb7ufuiy7eRT7tQkXzpE7yxGgUqZls0
O38hhDXrP3vx564v+szqV3sijJ8gVY9EaTEkXK4e4GCF6DlRAkUSQo9M6YwBOTbKvo9f51SKMG1u
9zuSbrUQMrscA86Vh55wTcMQa9JDw8O6RJ+2X4lyp5VGFN8mNV8oJsCWCg7Fghx0kd+1n3+VGyth
5L38GFKhA1x01aJRbcHqedb/tMW/FuE4Uut195KqyOrURi9IH+tp3X4BqBt0zOrhbzIoZK5e09b8
xz4oG6CJMRY2u/3j9JEW9Z6fIYt8fOWduECXm99x/DbbUaqRY9N3gbGk9cDnd6IuRAwFNb1eG5em
SyeWDz8TPSAAgvfiPuIGJOxbMsBvHG0aeU/Vx+OKkawEErq/X2R5lxsSsRM+kc9X0n7z7mVSUHqf
BDJfMfWZxeMJjO5cHSGXlrLx0LQB+6qos3ulU89KVIZQDMXlRFFH1Kq6fk/68hVkiu++C+fsmVIs
kji9cgGmgG8Zlr8NGglKBRIbYO2D3XhdfgZOrpsFSrF7DFZtaFErX0OSAfdFdlF8/tf9QoFowmJZ
MVQOqO0eM3vvbuQOdsw9ojtblwimRRaY4RjkK1/VI0taIGRD7U4hk7ar80881mvWJpGJvgJatuBf
e7+YSLr7FzhRpfnnGpcH79YRs+C/u2cOddT314OZ6OF941tYoOVIphyS6c2c8ZZZu3J8U6evHncS
RxfE6sxam2SqlxIW1YlZNAlSM1jIOFIg9/TKm7YKkldWUUwWy+hODV7JDfOxrMREi81orBG3URj+
ufWnvftKNbz7dZwPAT0QwiCDeWbF95KlStbBBfPe+pYDhL1wm0d1+Bob3Vy2lVgwYJ0g/tgm1+Ju
nLFIDqOWSaOBbABqm5APLDLdwQFgl4V4xzOAhY7vq8iLT0vXYphVyDJ5AvXW2wMaNYjGXoy62uk+
FsIPPHrLkoOWQ1ijXWqt46Lz3qFxc1kmV/WUI3wrvKQ0iFe7kKjf/ZsLx5zuEEzhxRKw6mIfHwH9
6pWuVFnJCvKxYK4XKrz8OwwIEmCsdFjn6qdUN/u4obciZq8i7fsH6OjjKT4WPMWd/JZfWz6MfkeV
c8pu5AtpjPuyvcjahUop1+aDzbe/lWzX8MS+QuyX7iWEyorP/sGsQ6c1qAPI8OuYqCGs0v3fxrpw
V6+4XsahRl/YqwqRIY8KtvjwX3jaBRNWMHtH0GMavD7WrxjoT0le/QVyJOEFfleT0tkVSVIursiF
MYumRXevbSJhpE6FD7BHWSMkj7zHn1mcAxWu8xuSjCAPa4X6xawYsX4YjOaKRW7aT4QsRYljLV63
W5qvhN3b403AsiihHWUABISCcVIBlDYMHv6idYJ4HC93z6ow0PxeifY2Jpo1Gh2aoPzJyNzgaEzd
SZXB8sO6GMnoqhiPyoqEVgjvfu9IGtAlcZMRhgBHLU0z4F6SI+FcN/10isT3Cayx4h8NUVI9qX64
j0BKrresODrB3LPzzKDXBozyB4IDtn4uG9fWmWniZm/41lcDoPxrbXAdQQMoawhJEA4eIY84hBA/
v01B4HXcIsSJUjB0fQpYIK43JPNqQ0JBqLXrVNPQqppvTdHHpS1yQQ5msrri1fqbHyeDosPBVIRx
jD+8fBibbcNxDf61ryhYk4D64bjVksqaWQHywpvD8UNW6cZ5Rsvv0HPHONe4aNRQwoDK9DafWwAG
E2gKvoY6fT9R9cIpW/CyxVJkRnMjaTXKGkQ6fgjH+hva7RIfO877Ikkf1Y4i/OqQRz+YaPCmI/mB
PAP5jmRwCynDbkE61cf5ZSo27ZoZFIzLWqM3VPOa4AzKMSGKCpqCG2624XiywVoIfJY8Ook00PWZ
khHToCkLwQSqqHgV3d14uTMJj+C1ZD1IQjIcmGKefdJVU1VL5gbzANot2DOXrrmnxXe0u5TzC48g
rEZDvM8Dhh8+6j5hWbh0XbuRXr7BhOHAZ3mRq2qKnMr0liF1BD2+NxAqINzem45fZ3a2qKqp/UoU
FW6t6GMXvrilWLLXbjDe1JN+UKSkmmluHcY7xYNMoS0LmC9ov0DuGjN3Si9+M1UxXCV/4tK+bwdL
u8/BSkeGmbkMqmPn7RHA+o+blKY5cYgi9VwRq6qEfPmBn/W2J4kF4+xCOHyN+fuP13JbOYwKDCHu
V+oysYjV7CG+Dix+geApG4uUUxxq/HRFrGTf4kXUJLmFFKf4i+68iTRgqwO2ImIoWl11eW2K2JGg
Fx/UpxMmSj2NiwgOWPGN8fBvVxA8rWDWZBAhIkYDsQ8ZDlCHkBeS3bybpZTNRdiwomw6p68mf8Kj
qtWsWXLTCFEckI5tmbOQS89sgvq5xRtbqRXcCZN5y0Z/ySu+Yb2VTPRU5E5d63Nzviv8evO/BsYS
Mxf+m1Jb3y1UYfqtVNtHvs7K62retYHJfELSD5DZhKwbaAtsbf+HB2FMrCuUYZ90LD59eoO6X3fA
gKQ2MJEhp0s8bj09JukTWUCGTc/vC4u5mSDsXuNFQ9BdZ5n7+ro56qT/x6LsWa/LVgQzfqBdFRAQ
qmcPnvlYuCmJZ3bvfMuAf/Exksh9u00ONJY/Hp+JWIOj7+lX9uJSXpb0Y4SqKQt3YSESW7uWxiz7
1XmlduZYnB/2ngL89nckqrDo4nhkKah7Z4g6++uoGu8LBSw43DnE1tZBOb04bD/b2LSgiDlcp5Mx
qQMGDC/QWMDqhD37Uneyd1fC65VEGIueZW5F2oIS0IkAiraiIMCs+xWfX6nyZZ13LtrWXACKlRwt
cHhU4+MSjOhM8AGBGtwojxj+kXJ41GHcsAzWxwG51wG9TxVQs977AAZBWt25JM44CR3v5bv08lnL
wDbjm/f8Y7Aw7+y1VtkG0GrqGmKhLjcPn1qfURIqHocPrzP1s38JIkAz0DeZgC3Yf/7rCPfqY871
4wgCRPXtxl4F5yxPMRPEp+VmCZvre22bIg6EUTUXJGG9BDpbM+W5MSI4k3pXIAsJ9jKxagw6TCq/
O6ld3fhh3y4EPVmJnq3LGmXp+zP17ArKNY7GkLSn7BN6nM6fA3UB6s5WUUiOePhxI6CVJQO2bGtx
AbtSwRK5QyzZ8DzOoKwzFAhxHlBzpZxu/IzZdL2lrbOdpZ/aRlujs7Z6W+43YaVPmDLkFSI4tTHr
u8GfCMW7Isq7gOeY2rkvpyg9UCqLqtmtsURNin+7pJye/7bh2y+3SJU9nOzyrdPRDvC+pSuKMUbT
AOWezQpVmdE/b5AcebI+PmrHBtFFtkA7DpLSRLi5LshfP11Oj8Y6C/huSCbUz8YxUyMnBLCHU3cT
TbGG7jzL2NSPEs7cM+aWYo5ogl2j/zWqHK2c0QZK7yqHBqwPcKl76zqO+iUzMO/jQLnqHFz+OZ+l
CPOWLBAfH52TdPOQ45gAPeJgOF5+29dx9D7u0sBP17Wgi2UAOD3maxwhFZdsvNCg61Q6lPk2FSan
1yI07EmsEe6FyrCnDI2LmFKjR9i2/pPgiy82/E+2o+1EIzUb64P3gRsxMFiQO4vTheupcdjVCCIw
KdzF2fmrxTEHEfBFcjftR9XxkjaBMIpwdadcNINTZ+TXzBIubpjIwKf36dsBVJ+U8rQ+Hs7kdkcI
Vx16psp07tbRZBSLa9C8JgvjYZxpe7GQ17hbrrzE9nbq+QLJDm5gsF09vYr303l9JVsB3yxGO6fj
260bsyo6mnp0T7JxmvoVEEwf+x+cmLFXMJE0930fdoyYeEvQQUZhBZQ9ygVIDe61yd+dSinSmPTH
zhUTq5nkomjKuu866CKKk7pPwMImjMOe6bgsZbns4jjLYhNZgpvB6JnDUugRQroF3DHbd+O4djNm
cEDbCgi/EPP1ZKILR23TK9HO3EhoBmzqMzglXXftXdydPUhZ4w0Ok7QoG10eB3rCM19lttI9IhSL
3KecdeLz32PkVs+qjsU8++0fZB9J/H1jKBMLxRflq+s5K+i7azNyLaxsF5Vdpk/+mG1tbHHem/BX
89t7quvrF3RXUtyri3rgbvSRo7iKrXkj0blxiA/Lk5EL+gXApaybVbFE8wo1YqiJx2mUJF+sunku
askPcf4lVA9RAvSRtYeb/JPa5hARRPPqVPCpW9F6QPhQf9RKrZDnwHpvALoHG5V1Rl96zOXmNpin
0qiRQS/VMfowhQ8GQm53nq4Kw8ZE7gK1nlKPBPeIvoUo
`pragma protect end_protected
