// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
TFlqdcbWMMECIdTVCWdE0GoLMjtlP23mGEJx2W+yr6MZMqgonhC2meria5r9xBCRSdSvlLZbvoxc
WfJ2kKgukg75BVGk11EWGrIfpEkX69eWlQEmxF3+2ErGLQqD4JeCr/6VF6H+2+3xqbqEv9gqd3cH
Le85qMsqRlrDV1ock6IL69kG9ynluOIKIjQlmvxFwS6o5BMeouCXExHTAsLRgvBvanNmEcGVVMDq
u0gqY0k1vc4u5vfqpvLpajkJuDmD+B9F8B1lZSniTiyvTot4Y9snNP3ZDAgBRbJt7H7M5EuTBtFL
GB+/OFVA2RFLNU2/k2FZGl+fo9JO8BNSdXrSJg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
CDJVB6Nm/9w5Y5pgPXF71xbczKwXC7WrpAhsG+hTsh0H8FWjR7wYh3+oKdS0Baj2kD+R1UYx+YAz
DeMmoDpAbY2w0sZqeit/ajR6uw4Us3eVj00XQMEOvugZsV5EJPkDpIJOpZX16E3dY6y1UI4/4cJz
QvlbBrBHMEjp6SpvCL6el8TCrGl6I5Escw3cuy9cSPedOa8SDwsgUKm/v0cTFxgoRZ+mw474oqwz
ybna/5G/QjaG8I8Tf0WRMlORoRGKLw6CKo5w4fV/V242RPjW4mcJiQs1I8WpVG8xqq9YOcJV+h+J
1//tDHVaufFwspxrQqUbnrQgikRI+ggeWblVCk4HTYTAU4xW6bQk1vl0n52BJajqKArOxt0sbCEH
2jbgV+aokWlZnHfHEc4w6tBDWptjCNsPNqktPcK9CAIrYHAz0DyXof53/98wG/NFQPBOri/zLvbQ
iaSCxRHfG4PvsCE4zAEMIl9qmRhFuGMqBlGg+03ib9UEYYrPZ/HG+C9h1P7Wf1c/kuJOiEz4l6tC
AFAIZ77fbDwjVWSt8qW9AVpA6wwGyCP3cJ3IWOpZxJqoDR5f2y4987NGtyXzD4TiBCFnapJsk4uL
IEDZMFlmhObkAPPpf+sn2FjiAI73WmOEn678U9RTlh9nftspXgLgfgCKwwjzzRiXvoQR4Ad27sYA
5ubLbcZUbPzP43kGfDCWSM4C3MnXi2nJ6RoaY2fFX4T4wxEZezUVvQsDpf1xr8N3heQBcKvzL8qb
6nlPuLzsfAuMYPP6y6m6rvivJgy5hmZZsqn9YiJmhEZTd7dQLrRWXbVSivf7DIrmZdTVR1mFKFEN
JYM1ByowQ+I2NZKeTBqMiDM2MCPNyBjOwuNthjJkLrQmbr6MXei7q3uBNKJz26uZkrWeSVLtH0pP
aWiPJDthHkMHbKTGJEpJlvJUnDMxj7bZnBTIHV5DDRtweZs/n/74JViUKkg99gOMW9pvrRffog98
Qv5GB9kp4xtrPOK7gitbJ8goMobk50VMI9zUqDlpt2uAbrXoEw5zXv1onspfztIR8HGZDvAYkgGF
rdL5AX2lYh6HnohkijVOpVUMWXLBUiRU+7AUMUqzQRWRIob1TiLlAXnhA1TFCO4c4RaDLfIx6qdm
9cSyOp0sto6RJ7avRK1lbEhWTIwStBvb85hVFmdeKc+AqXnC3rNM4/xT1iPT6f0CAlD5eHqSSd1C
MjPBpm669wpAR44vEFxNqMaa65VYnvjSWdlY3OJl2p7Fv2beqiVaRBdsS+kjqnFT6fukQSLpehyD
8yGiFqIZIn7pe1ZHVi6MVekYokQz8AuQEKfV4NUc9FAzAvpAWKo8nESivuf3VPRSrbU0Q4IeplbB
Vl9GllKFqKWcI5Iuo8ANg+Buqw5FfV5UGhwWntRJtD1IprNm3Sepn+uA+ogx1bWvUpDKZOhb4Kiv
uzXY25njb9acznu4AENszuR+5/ltsfsxaObzSa6mucPZV7m8ebcdiiRvgNNZR/4jrPH8olq//prR
P1Nqq2AvmgvcRHf1b+kUVTHJOi6GnSjGidfgVm5pJ8YeLErN7naAbRdxN/YPipS+wNMaRS+XpIbm
Z78yU3MTt9vGVA0UumFaBrMpp5bNu/cvqjhd69AtDqrEMNtfSgPl63QRLsRlCZSP+cLGnNSuG2NW
l4+mfhZ0uOTs3YAjjft2hN54uV0ogGCr7cngv6SBranj8NsQWmrtYkp/zb0O9nFNAhS9J6gWFMWP
NmeUNAXh/MRyLZjl7M1Z40cBMazM9kXktjqf/IAxUSSwy2w+DibE+qshBt5DA8FRAtqlvM5DCi51
qIDnDfKhglFmdhMlPrm2iikl3MCo3FRVmo286hM81xedoAOfQjVi2jWy5WS3OyxPlYm9vQ2VqF8H
jrjkFwW7ZbqeC+rSNzgwVIVwuAV9Np6vIU1cVXNulpKgPUQQEHUeLf9T6sH6TUmowDN+AfeF8d66
2FlqyU0GuM5LHeiHurF9qY0vFgIf2H/Kx26fUB5TjXHr1hRZ96A0Ej1FIcQpOL2AXKrj2xG9Y+36
wezhFBqsv0ZmXN9mErf2HvZ9XMCTeGeswIkNKLUBDCnSuOYGfzHPiHxfKXtTdCqRHT359Je1t9O6
eoPZJGoyrpdyPlcImXmCr/gMi+p/PV3r34YVmPdiReHvLn1+BSd8yWBSVJH91AZ/+C34LB+15v2Z
wNShDrOQVlnhj/iAZs/ajTU3ukTsNfcqW2cnGfQC7ESTsMW1SvgkACgxj3C3abUmEROd6e+XfFD+
2JYv3BjHE/DJNZChyXJTEzF53HcwRM8ytmu+L0+futiQgZhWr4G0NE3TC9TQI8Zofea8qTd4Cdtv
Rc8G8S6II6bbJhk7yLB7Hew6vdW0Ox4k2QR6PYDQUj2KhYCsCx+ZEpfgoUPxjb6dYonClzp2QqB0
jikbz76Tg2eNDYmXyMN9bYJaE4sgWojvDb8TqTzYkl136J7q3+2TJ/LOXxqCxApAZ286IIbx5N13
d06s1/EWuuC/oJ6qc7GKw20WbE0T1Zmk+VqDf2/brlWlAU0iaSDUVj16hYicChI+rXfDMdB23oHw
aUpIP5MfxFAXOhkFzNotMZyvkBS6a5l2YegjrbFrD22AFOxrylMPmerEw2VOVCjDxXmJX3PGUlr4
KLlMPAyKN/OyIsgX7tT4eo3xovvkghqYCyJrfIDR5X5lXMk9x9lsCtt1mBXSeeSBW1NwDkGhmOvO
Eop6sjtGX7hOz2xtuR2FWwkDfm/fCc+aEh+4Yzu440t3fWcovOr4ZAEk5appv/3j0QroabKHRQa6
JGu1VTW18lN9lEFzEhUunt0uWtdRn9G8ltJ2VADc91xmecb3naYi62HiAEVXy0FQFRLywDqnHFaP
K983TlPKg4FH1D7o+WB+EjoRi4fU5q0Efl7nMxRUCcmXZ9BlZjmZovafLDcL9TuFQ12OrGSgligT
kKWIGj8VOKxn9lEypwNicPnvGgOWUj5756IT/WjNJe+c5rAs1xaEyAPHictvbilzp5OTGvoyRNq3
/dvZOeyNndk0wych030j7mR6aA0hoR64J4Cv7JY9ock7FTK3Tvtesda8OlHz71nsBjmcrGds4LrR
vm4aKCOPaUvs+GA/DfTY2OtjWrF4uBv0HpEJGThjWyQFcNJNWcBk56sk/VshhD5OQ3IqgUAjy3x/
aLswDiv2lA9iKcHqxEER6mMl8mbG988uir3OviHUHahE78asPKo0JmNVImpgzTWJ5oHQe+5WkqSg
gRLakYTkTAeyo6fiWGbTbtGrQgjh7YEZkf3bh/PTTojJINV7b0WuWdgDECymU/hxNazxy+q4fWkZ
xttIXobqojQxrS8lbixhGjUeYdhJgvlm4luWavWkDFQqFcEJVi8zE/JTnrVzsX0edsT2/200DJyH
NHK+2YGeM4bdQODFgRHgrfLAe2B+4hk50oEjqP//FsGDJuCEJ1zM3JdcLDMuF7dFUaiATGMZ4DZn
K+TAuRiBHntHpBnn9Y/nUBDfwvgG21kYx3FM5O+TdhT8nvXCX66nxeqDtI9TJlYjpIqieTWIeXfD
tk4AYdH7FRmZjeJuyl0dqM+JAFYUx9bH4dY66F+LPI3KWUykeJ28QzOdxqped6B1s8Z5l8QscKw9
iZjKh+vKvm4ISPiWoWPhm+2NnnzYmFp6Wl3cfJ+AhcwWrXo7EyGfsaMG+DE88p/skskctr+fx9Xp
eL1xANcgQ1N2p+YAvOT44rU5TNDKLiWW9H2uKDsMdBIkYlG2XDyQbmBYRcuLXKI4dc2E2MsvP/Z1
gaRE3jJKtNqA5gOtUU2wwqB3UVekPEueaa3J5XUyqjZ/rvwq6RHf3ixvEkHyCftjf27YOXFpCRih
ke8qCxHpKAm0pmvet4+bwB8HbNm8vuzVkf3fi533sGxbNfayTNsgs9zZuE+meIuswz1uhbYgwS7h
r5LBOCj01bmbWhiXZaDDtJGFTN72qEXkz9f9xpNljUCY0lneXBjVy4lR+61XZZzyBDkyJuhdlagG
kVBpFQcx8f54aV4vag3zSIqJdGvL/6dPkV4vfdR9HWhRYGSCcZGAsif9zJv/zkmlThyIHebDFx2W
Q2HwyPDjhZA9kUS+SVR4h5T3zBGL/gPBnY8tuoaa9hIyjqzwelscQzvkvSf7X+12CP6hI35ZYUS2
nl1bvyhlmqOGZmnrpl8idtnWa8P+9TIJYfBCHLrOoB3nE0llRYeq0joXluREdMxFczK7FX+g8gsB
4i+r6IE4AxOFQU7cfT27sqEjyXwGywlA4/G45rQ6G7WSpHhY1D8gl7OHCWSYCIkRMcgxcE0tHzzm
qHZCQfu7y6sgeCeUTGiMgm1wuuKD1lGYvBKK9aILDCF2H6FD+qUkNTUK2SePsWmhcJGPbPIJfR59
4Dqix3yJYxo9f3b0kZvZLg1Tugc7+5g5y3BpJHR9nyAdvk8wveMUS0ccUhEKGnCBzPl0vGIHNLP0
0xf0cmdoK7w10S8Dn5HADFKD1Oku+sF2M7IopTiF2CC3+SeWVQGZGpbEPnyzFTUJCdNiUL6mLwgn
lpeKfgvSt1fwqsHWK7twmxb/yDVKIBYCqSnuowv4fJ8g0YOj/d5PTMScejr5hXN9rFSbmmhjTSCd
Bfcz811HYN31bugZsPlES6UxbuAKLXA+0lG/v7WFTXskjrm3+H0W6O1WXUWRp6V1ady2/vsy04o9
TQRoE6XD6ZkwR+DyTg2oC2Z6Z+Tq9W7odb1o7/MT9mrHKhsSt8s+630OAwqOhRItwd5gM/qLQMDn
+tzELrSjKYascXCdvMSiHL0dQA58KkOfVzDnRAwXNqWhf1rmChU1iDwByWKFxC6zcchHYAF4qQHX
Yr6vlC6tERxA48DVyfUa8QKyFCULWRh6f5vLSAEUxIjxMomNIkOHHf6LXgqcuy4yUsV+oX5ltn7W
WrE2nOh9MQV9dccKa8Nj1ADU0HGw2OhS1gzSvEwjzyej4Gwpj9MQpvigp+l9poPlxKXnN9FmEi3d
yGvKg/Vq5FipVnOOZpmiVHhNFmSiMHUqEtn7bQfJn5qmoJCr2CIJBl08UAf6qFAEB/vdNSESJmQx
prpSdb1kjc6zk4CuD1jxHARyGI6SYCeG8YEX2M7Z0ttK+TktbpI4nSGfYHazZglaG3ruDykvGSh0
UhEtmlnpqcihDjd3Cg5IdG2uJb1A7UKhpNb02+1iAnKg7pXv9ZhfWwk2LywW9q55YwrEpa0+FnPY
q7CERQD/k0mjKVtw+UoZct82ugIMzvNBsvIkywMfWwE9u4kockbDYnRFbpRstVJ9zcXp8LPutBQN
y7mnsrwAoP7tNVssebeySOSz8d25Xw3Tblov+hJrje0ViCrby00NIYNRtR5BwbulJZ9RCGbC8kWO
abh4ZCh6Op4zfijMz4NxIBfyr7RuogHb+BHQqdZMzs9QNGQImWTLGnJNswEniAbzIzcaPPpJ6OIa
/aJkGnY4fJzJyxv6qd8jO5JGrd0cYp5ruMpR4M7VZOT/l/73Oy3iOVXjnu7bevTwXhoyzyYlRrzX
BO4t5TidnOYzu4GEVguXQy2rH2AJA+cuVqM1ssWRDtFgRIlqhyaNiGTYj4I73Hr6gZbP6XCJBzKO
E6o/HaaCd7ErLXFAFxQA40MerZz46AI0LqFYyUBW8cQfsew0gAKaP2hD1MWiws5hXlBvfCTb4B+B
hsx9DTTO/DlWrGdhI9ep5jPlj6T0xLvG1k74amOZiKmzVRKM/gwA9Q0CNeIEGFVULesm95mgI5do
cG4HLXvJmG3lwYfoGXiyv9rsPmdXpmDxlSpsJkJvXd/2WtFjnc9pEpzgzFKdPZ2zKsy1DAT4yrJI
ARPTmUT8kiqs1fZCir2MmXifWYpnVBr/2CclZW3rCcgOQzUPKagV6JhZgMT7cvvu5GynFjIVjz4v
4rz0hQBXkrPqgfMtSWAwyffV1CjU6cJnAEGBjL1+QZpqxFKrsNrxrRRXzI7tsQk/Z9LkVeTTAid5
JoV+DCtDFdMeCl3L/Mwt7dyt0SmKIq+WrTp/ftPZOcN6DrsuhQqT3L+JFuaZe7aAeRomSxJ2gI3A
M5BrUHB5QA6LHnmBxxaHCdSDriBttlkCDkrdhpTxO0sWhOZB4i5KcLChqJ2L21foIeyIwNhyuDtE
KwigxyjVSVGqMs52C0/ZGcqd2sDIaVxVvsG3CZMfaaD2D2rVxhx/ZOSMGnRVhReJ0Yww9tq5uQv1
Lnl8nXB8s8Xv5ObV3e8ZVcNlaDDofSUNLnK/ZgQoLAALtelJkNCTCx9B1iGbzI/cnc4Z5TEZijgR
iYfGh4XegDTR/8kHIJcJPG2PURrBFQD9DqGMp0h4GDYmGpxAMDwZniaeJOhdlnGh9Si9TCjGpmMo
tvnVcx0v6gt4W/BPF78tWcpY2b5H45Tw7wpShmJ7hL9G27fPY1SiDX40aPu9qagZCpoxKPolbMyA
thXW7OpXoyQsoE+XymcLNes4KWq7u8RlqSciGV8t5HduaskGCUyhOW7kUD83BfXGX/lADGd+0j49
8A8d+Fh4FQLwUBbQHuzM/qB6LR+f5ah3fKDTRTrL6v4fEePzo4Bg3uGDswLsjWTfpsVCFVJVmYk7
ecOKQKZhkodJSzGPSsYvNd0QrwogKZElvsB7Xy1VK+iA5L1w62fYpODys4/Z7x9O/jBYTTkyyuFJ
2U/QPQ6kQR1SPkaBMx+dur6OkYmMxRvLfAIL9vRbp3GaXwJOABB/bYjtGf8v1NV6w487hi79KSo9
VrbJcYdCWF0YeNqdYWiH547P6H/IPgnt+Jqm1Bbk+TAp1KDvaxbCozHoXt5RGR0cAdaWVyQ2YZFi
i5P3HlCXBYLge85wnVdaGSKqaA7Wxy2RRMphnjY9I9ew2KYWKkuFZ8IN6yvMzFdxkLPgrlHlURGc
flgN6eUuDLW5dWvhndB+DtjgI6MvHCiY1Q6ZY7frFgG7DjBIhCn2XXDzFXKibZiuZDZE33v2utf2
y6EkivNZDsT4K9cLV9EAZHtFXS18mr1KYyEurrga4ZMKpqVpSTdGGPEzDlxaW/k+F3cN6+1G+N9q
3F3gxgM52/9jBW+jXlF8kqJ6LTff2BDtZ3Hb25GPC4ymIBqVeD/uF5rvVl/muofYIMNFBg9yqqb4
rI9BglM+CYOKgmS+b3Ni2JOSI9kfy8IcH99rVMsRtXaBe2eRiLtVwsqIX/kd9+jsxiHuM9HGx3wk
wsUWjidus8y656q4dI8+E3mtSlA5MZWdBW/VfoYAapWIr+D3oHgVG5qXYRD6++vMWbYWBcifcIR2
jEBTyamXvGkrUQt/axpAQnuQ+r2Dsyk2xFmDqjfW53bUdRpgSvFUIhda5gR/h+PSY/vcpXZEQSxC
bLSCIgvSH6+N1kkwZnhu6UbNuLCnmVln7IXzF6bsRfQ1r0H5COxcoZ1Ozt01Bq9MMBXYsdB3gnkv
VWoM3Dp913azFzINZWLidhnELKsczbq7jbFwBA0HtaAqTksiW5tmVASuUK+ezekbMW0Gi4ozdBzc
cJSvu/UIY/qPTD35Ej0b5IKVatnBF7HUhEfzNoh6rUdKRMWVLFAcpsgg/7sQntDZMVlYpQfL3Iiv
YuZrQTs5D6z/h64FkZF0nCn3O/tQZrg1LVSpENocaMjE0wrloQbUe4ip5aXwfSdqGwdP6B4NBTL4
GUA8Jr3EU85lJXM6806d3iYw7Tx480OFRZooxZ6VDkCFahkMia3hn3KWI43egZL6lEpFyOBSYS0W
vz4ibomR2QYwIwR8JIycw0L0dh8XOg7TiuzngMJlpS8uVr/OyHl35f23IRT0CTPYHgVM2l1rpYTT
tXwCoTttPKUZ+6H0FNX+Ybm+iYqGOMCOByoKfqjCV+t4wy6KjoDu5PDn7eT4rtbqHuUdp9Sn37OI
9fEDaae7sW9AYufM3Zotd1GCpqUuxopA3HnGRfSv5M3pDOC4XvJ7RYtbEkAU/xkXnQhjexce3MyI
hA2JL6u8/awevlppK4Uy4UiUxcoUdg1gW8j4PPOQ30oeFFK/J5R34q7bDwcF/ZM+4ZBNQm9NpP82
+JvMEujwETLAmm1qExBJHjVBy9v+cRQDAlCXKqWq//tWdXCkx3NOUb3JoFe706IAodH0OeGC0AjK
osE+NcJIyVpvkaymfUlRtdrmqQ5ynZX0GCHSjfrH0a35xo7LU1D5UXfwkEeM7OpeGlCVK2+f6RgW
Iwy1bmpO5/rpmr7MksjiqASXLRL391aROD8LEbqSHrgO/08AoUJFBIChB5QxrEGWfFKQ4osZUeCx
I/WQg9hQiqwA6fxd3hVZGwBJ1Hj50fDwnp9ZEQnjmTAhgkLHC4rG5iMr/B+QcaLQYmSBNwtmfj2H
XOst0iUh13k1IBXyS/EWvmT/ryBxDI1zJs+UdTzyWqnm0KI2dnPrDa/m4nNllT5UgJbSuyrXii1Q
vHhTW2k1UZ0jz/hcWAkHx4LpepXlxZ9QDbnm6NX4nGNPnZlnK3exphOmn8eMpQ/n1rUNjcF+9Ngr
t8TuLBynbsKwMH7UnuM8xIRbajDdXzJ6NXNJ/3nZpQdsmI7TMbq1CUUBW+TzALfCdRvkQ5eSa+Yv
Qb3vq72UIxiwiesvZNWl99dML3jR2Z6s9mFv5Pwip6GQJEenYyLEfTLTRm+TiTqn5s9x+ND/nSk4
HOIjpuG7XxNi7jMH1CbGsACZ3wDQdTEcaxRJz0aD8ovaK5k49vvjerthde4Fcrdieblnw2m+8AMr
lk1Z79h9w6otu04WhJFIALRlA+EsX5Y2evG8quB1v32q7CXcz/gJQZYid2YkywlnL5ouDnxqi59V
ZrhaCYnHX2FNljyi5B7hfJCqZeFT7HAH0t2e098GRpyOvaZnFXCEJBOZrzMSmpvDKQnOwJ/TZbJ0
eAVIrTQDGniIx1aZwcUAWlK0CcV2ECYHgr5ZQrXoSiH2nDL5/GmIeEkEupJ6a0TbkTip8u7p5sBo
I0JDTlzOis6AyX9ba5TRIDUMijJD/UwG0JtMHorFA/a+a0fdxNEykHkR4DifHp4F20uxrBCyMy/l
EJ8OMiSApvb/YG5leKWWM7no5d6nkSahhDhRBtD8aOjmCQ8A2d0M1LJcPUEP1yaUa0ve11dEUuBk
wVPPFeqR3vViae6v3fc2CpYy5qNiTI+ZDxLUAooUDyKvekYFmn2sqt+9L4cmmem0JS1l910087d9
qTRwHHDZqevwkyTXICQqs0q6R+H9fcFJaMgNNt5IPTYn5bT8FgXqnOCdPW6tQhm5F4hH35sR/t7R
4K24Lux8OroI9p9S/3dp6lCxHio6j6oiW+Y2HoIh3+XD3oIrSVBGSzPulJZqn7BxI2XGYg/9D2JW
AQ/19iIggmIGR5Gq12TMzSK+qIgxfjE2nw1TgrcoQSMetZAorTbTQK3+5gX3H+/V5vSJyUj/fP7x
t214iRAGATUCCcdhsZFtq+K2rHUW7ngqOZ0HZP4AtUrvKK7pQjLzuzv1J+vWZe10J+JvGMNVDr0M
XxVoBbdeNvxAWS/03fBltTM/D/fmyVyf6kUUaaS8SDIZWM8Y0mEIK/jSlPVDkufgUTCP0/a80yEw
O5THankOclnJnfK6a4Lc/56WN5N03rVhPmti7kqOFUQCuvVhGfePgtA78lx49rgIn8jF1bqZot9g
vXiti1aicIuSlqB7CVDxytubqptwT+eZJUqcA+qkdDiH7+oyzbbjH7RtJm+f4cxnk01hDmRE5a4s
Mes+Fy5dvaTCvmJKWy9vVYqs8kBEp0NMxBPEJ407gYxSZKQTcqIPlbH273c6cIKvEiAN1iPNLe5P
nDAeY3vbmv6QeB/XG3norRuR+G2U3fWSDatxYyzO6+8tXmCHtyl8lv6c2kn+E7xkFMWulz2q0cKi
XJKFz2FhV3xTEAilI4wUgnHqaLUBc8/ha3z3k1psIbAIMtf3BKJ0odHyW7pnr3wutH/th16Owqnw
JmMsrvAf3kH4UJ2haDUBtGhKb4U8K31SW97qwnwTP3ON/wQtSyUGUdzCL2s/GyRStfPW2eZmIJWw
nmnPqDqKmkXCUi67E3QT77eV5ZEVVIscff2a4rHlg0sgZsJI+ZNeVozndrPB1UW8pEQiHMFf5oDM
BAkDjveltrMoIuLew2BoalEDBXOx1t5AjNM9qFMbVbGg4M/X8RDvI7Q0LJUhOAhu38eJrouqi5W5
/XZmNpvpgznokshte89H/sn7kLEuqnncN2WsQGmCXHREpbQ/tNA8MbZj+BKbhat9O7d33+owlwbM
Gw4fCQOzQuTaeU1Ypc+R9ER+2u+fQImfkWCYGWLUShbXbq8+ltkz3Eh2OhD7e92iNpsy9Er+yJRl
M+rOMiS85uaXleIx1cjEeyiD1f7WVi3desoKXCNmyDK3XcTuYqNyLQLyCAw9VQ7sZi8Lu4bPIOPK
mfuS8csKEPPIkd9wuSIvuf4YJNFLMuKVtB75AhG7edNxIecduZmAUU/Sags15axFV6u2l5tXhHg2
pxVTh821vV5PkKYahzefTeLXQlXEQxAjj8SxrWf+9tsr68lGJzZgkguOBYr+VwymFDR/x0KZ1x/y
tQFJGZIp127HnOYXUTdiXjkRlsa0JXjTxw5BQGysnoUW5pqV214kwmOFgj3G7r4Uel2Opg9nWoby
BsF+Fij8n/ZjNfTYXjcurPUTZ4v2l0hn2324WCUQUlViCNoYPRJ+atfcHRVoUmYuDalpo/9Hsa9v
4f3JUmevndmrIU+ALJTmJ6yPU8sxwOB2yu8bYfmy51xwuc6SZF98yG2XYmPoNlyUhlE8RaaOIaB3
xRBMzT3dF3YjM6rbuamXDjqsxWUrDcNFgxAodmyObnrnjvGHvZjxrzlAtPZEqQB9s39oIcOLWMKj
dqey6vFKMyj7fEIFEA9plfbjIb+edCmlPqsXKgv3t+5HLf8y+ImhulKDTwJU9SWWnjYm0l1ZDbbo
vh2IZK/P4ZAU5hyrpP3K5Hxk3Zt1ZrryplA+EA+AM9bEnDM9INnI6sBi4UMrqVfh6tk+/W2ES39O
dab/QbkV0TGwcUKqVbKCNT9WNw0xs1VWuF+wNfcFO1M/BYlamspKHh4u3QnjYYNvR6gmtpL9gzfQ
6Ir49hnRJa6KOmTrQ55OFoO0syTkTW2oITVfmdUTma5th+ea+CCBsxZ0N1/mabM//5UDnq/NIBnF
VChHTDvAz9xHx4443B+zlIE2nqV/0qHAutMFPoDHffe3ZUjJOFH1du+b4UU6P+dz3pAIja/EdhA1
63PYsWQtOVYHnVbgeR4yS4AScj4tYeeHcQ2lgA26zjSmrLRk341V34mwnB7/F8BlMbL9PEcH6Emm
jlcWVTdLru+P0ohErtnjj3gnEVEtmeLTuxIkCin/Dm/Wb09CLTCSgbu0++eJP3Ic3+dfdeaiWB9M
qIwPXt5OCmbAhSQs0t+L2mLI37x7QKySrW7HGz8ChJ7oyAtcc9m9HiaCwBVbUw2xXc0j5qloS4MW
ngE6EJWCE4pYJwTwONqyrz3bU2FH/qVr/wR5HATRL+ObshXd9bqdiHjG12Jn6zX7G3f0DLCUiul+
npiC+XIir4QORnI70O0hjy3nqOJD6uDc0LCGQxsKjbZRFAeC0RSK9ziBys2kqVbDYDiNpb7Ht3CM
LiI1Mh/74Hr7FID8QrcK8cWQOEcbUJRpfbqG2bIj061lkbaPkGNT3REnrmMVR1/+R2kFsoingwkk
oPfOfuZtPISGpAKxiiRtPPBZgSYA/KmxfirFfejlKV9vKVEJl70hBlWNJdhOqSdHdgVCR4Bksj3p
fFVXWbrWHalE977HRdALuilfXddjQjB/bNZfcJquRT1m7q87O3uqdgKZJccOT5TH5SGzy+f01wL4
T1YjO6cw1+fbTvk+0hnbJF3ZTzYH09e5tD+QXYhMzfttEflfV8B9BqrG2d+rFaIamt1L77v5Whx4
6man54YjhjohMBtU0vBsjhmHBtuv4+6R4FS4ghpcbS2FXwwmoEMsRwckBKS2I2W7/2p4RMUidVIT
cu9uGl3IoZzf52Q8JdS4HAJcuJ+ju5W2Ln5+bQsDPIcnXy5fizqKCeo3w5dAm2+H2SFcrWfYCK9h
IUBblCvWFBKG6xavsAx+yaXvrWs6AcYlWBnCDnwVK+pYQPxV5KqmP2pvC+0TW39aGYlEUR5dtY/S
b2CG1BxNCirHjMPA6whl3SBo6pVQVtjd8yw+lzBIMTWULuU+uYQtoTwb7zNeyZcxNXJtYegfNKRH
M7KsVqjx/+q5OlipjNDv+tT9DWnZWhDOH0y1PoYHcTyz7XztQQkyAGhF5RO5Iq/bjdSD21z4JJ7c
jsXyyBDf5k47iyxCiUcc9bgJ/jJc8RD325JYK0yMtVlngiTJ7HIEGbj2kUwtfU5Mz4cCDukiFttL
Dz0Wujo54UxHPMYlA/KDnbzX46J0m9qDoiJp6y/9PaECXPIaAWHQDqYyoV5+G5dU4Qqg82fkf1rx
GJ7WGhPP9OeNSMafwgU2Q0tMPuAfQXYjrKC+WV3K7b9hy3FeXkDjc1Q6B3y/Pvnn6TWOBT8222R9
cF1r11j39H+PS4sLN8+vul4qrqH+4TyuaA+m8jKiOgIlEoNOoscxC69afaeJGSvH2PlQsA6Zn0E6
SXDuF8aD05olkSgvlTHM3f7+3b4dASCr7pNTk3GCetgcrhz2KOPG1cDZFSjE2/GV/M8zPjDUkLo/
MnUe3q9Bl/B00uOqfhZJZCtwC3iuZuDDif30efmTl2RjXg4koT70ho3fOyNAB7Bj4PU0Ilrue0x4
Y/oiIKHbdYlA9SVpwxdnucIQSpuwR6hx5vDF8cUSTcedjq/Hg6erkTbnjRPBsoF3Y42Ozys6vVS7
YBbT7mHkB7DoHVoj/brDsq37loMLuniltUevo7Ow7B2l9qjgiN5JNsFnqLUj1Bf15aEwQrYiY53X
YzsdY88QLNa70GTWJeYPntoE8J7aJQ0yfTMlE9k/zDUmdTnQsXxSwva5VNMmfAIcFa9fLOKAOZ2i
9suSNifpAD+S6+DvUDwpi3EvZXVQFq6XUkW4510YkB9yAX+pICe0w+58Zibh8mDNM7OY4kCUR/iI
jcLnD9SQft0YSSS8MIh457i52la+gPfSq2p44ZMU4oaAWWl0enf8PNdyRSAtA8UL8LwfCDwMGFBU
l6CZHyCTuikuNe18e52fm//BTyfimREcaFW076rBF8VbmX3KuclTJs51UdW50v4dl7jINxJ9Ukaf
AUT9OGJqHCS1xQVN6O76PrZFOFEN4420YIy5VoSV0y57FTFkxYuUDuV5lAzZlDkTtKdDAPAGsCNI
3I+oRwrpKMdKe70LPzv9xdOjGioh62XXxB/z1RMrbYWK8ScBllmPgLZO4k9k1ZiF3TTDR6NazXUx
XddkMJmveo7HgNPlrl/RJk0Bbdb/ThaFn9WWPzjMXN/4nhNmXvdU26mEibHg8RQiNEKd1wEwJp2m
BFaeuv0AqjTlz9HICKxAi2Ax2IVcC3UWnvT0MHPItKGqVmgZX48DHoP1AsPO+1H+XQhIz7Am/2tF
5CghZfEfSz78jPA+0uVeAlAl6Ftcm130kGEo4P85kBhTSq/jG9+/JUkPplTTUVzLoBVHZXoP1X4p
HLVqsbh7xfrcZcjV4O7ON0Af2K70V1JK9ErpbkF7QKuqdxF7aUXutSQmAFuHBSfpVrDhsCyf7qWn
gqAP2oa5etfGvsBXDylVqPccq6//HCmkhNzLLB1CUGvrCZ7JVfvHWMpB9NWDa0I39cKEtjY25xRL
zhcz9c7tqA5tMOMooK9F/tZ5OZIPlVgfp60W01L2xjMBebC3+JiU2KH72PbPKBYMEInzzp3+u2E3
6G8us4Ur/ZXXCmUg3s7Z5ttY/5ryhtzYw+kHTi2zNnCzl3WaLaNLgpm1p3TufhIqsadaWhoia5o+
Oc9KQzMnBzCtPE2Hxt2WgsY5cX8H3EIsU/BvDzmOCnacI9g5I8P5jMi3Liqi7URqqDM0eZ3QH8mP
vME4rQ2sGupiqp5j4LGfcUbsJsMUvijx3VnU8yEheGHtJzdeQLeiQFNsw7N9lqpi9rUzTun7ZWSx
8zsI1mjea+QfOfHZETUC0rtvp1JNMsVgQD2LgLGXxIao2k5YiqFeoPH5djfRsmi80FEwqm7+v33P
0X6g6klLmhV9RTq0SbVyCRR9XAC5wimuqTdX1FKLGpmOeTDwwQrvJFHiMwCjasnEl9Yc1t0dPlJ7
VKYLCc7AZBRz1HnzOCszEUnYSpC46VdGj1X7bokrs/3IPcSj4uho2WlPgCOd/cEIxRTonllC6lQE
9k5rlM4Y7Y36LQqAtdj6Q2t340OLdft2JCC1HzgZ3smhhsudRIwmAb+gtNsg9OMOZ3eVFHM0UIFi
2i8nhq+rbJ8COC+z6RmuQU2twkK1fVEW7p6vaOf7cGsswD96S4aBXn2WOxZZi07FtNTw45VL8+28
NpBF+sE5Dalvna6G1NdIZE5tMJDtCBQT3JtHpcq47eovQ3dWMnVY4JHbM8oZkqlRaZiU5VpKaLhk
KZOfVxwUdRL33ZTygVmiZf7McKo2DQyEknHbcJw5t74ENy1BziO5wWb/TUEzEXhalIxrEY6xB3v8
dOM74NUuIcXZuOenGfMQZBfJKG9lGoVX6XFA6R2pCQvkqDm97g1dzro0TnzhxR8RsN1rgU6c7aIt
Qh0yKHaj6qeXUNN1en+UulWQ7Xi69nPMgnCt+p9Gt0Sr6gk4zlia+VRiMyCIsjt8YsjvzVzXLqxs
NxbqepI1DQmiAXXjonP/fPEzTLWVGjVStHI4VuZxhTYeNK+ggle5WEoZECLGauRSms1lr/R0X0hP
3VOw7AZpCCswL8o6hsA+ltanoNyMbfU7wj5KD/++35czm1gwFPxxmferTcjZRRqQv64kLSPZz4Hb
E+guclzMq/rZff9eAK2Dgks/3EAKcncJBTHCnlYGphThqKp51xI0dr8B2uUUL/07KxeOCmXxQ4RH
DVKe9/uyQfU6/qGxCpmm6O36trKSzlXSu0BaB0u+FyhqOobANBdseNkSWWpGvmKJrp0HiLd9enNc
nQKUAejmXaqUBD3dnjsI0e3EK0MV8dL+QPQM7XgCRddnIccLjZw+atrpjLdltJkZHskBe9Zjx1Hv
voo+nz26P94UfZvPv6X197EpTKkMXmeA7EA0tyPQQ6xW0vgQBIQ9QyZ2G2ut4w2EOmvEEsUIPux2
DYAXbtj3AV1SzNblRnZk81eCX7RlOBPXC9DiR38rQxQStwg5cJHo/CnVnTJVqRhBDvoODNRa/Xs8
ziLrY01a+Mk6bz2P8ZSPs+l6+AwtF4FEpqRB8NRTTXklqM11/j/1SqVWqVTZ3QcDFmt0MqkTkEif
ZDfloKqbU/QYiIygY2vcN4SfWR7KVnDCnvwprzUm/Rdqia2/5AXlVoDa2UvyvJlXpy90pDLRjYO6
JAaKfDsCT28mCS83yQv97GupLVzTFUqi9ICVODWK3FUZHntkxvRE+CQSLMCiw0/vAmMl1nMuc8Fq
enIJrdQPP5iR7/jQqJxFB+Jj6bJnsfmb+FCL/FlqUfzM7rTgfK2uVflwjwwIZp3iouekUzxXc7fg
/72+VI6p7EfyNJFMKmG6pz0XM6FcIwxSOHVtUFd0WyeMFcsdDpm+p4CZwt//CSVjWTVo420zJbVa
19mHCojjXWnmIv9xSqHJeKIe7aEW+wDAqtulvPayYxUmCDgr85CzpsdCk0yRgvn6MyvfnRmI6/gQ
p3uv2EXEckc06cGjVoMphY10lPr8FW+Q6byZrFGh9upcM5tG68+BDuQlKQw3v5oduC2VrIxzfQ6v
gx5XaHyUWctPNqEuZpbaIsqqjF8LYTG2QIzLMvEvyzJan0+yGFb4UVW/DEC/1y+PQyfEabWh/XMt
VER8XvluQDX4rKlH4Rj0cmPgyPljcA23hbi0VNG33IfhraPksCswqxafyN8OqDWFdAbgyqDvGMqd
tfFzpEJP4/n7zBnru/ETTOQmEo47AjRC7a1L6RapfKqKZgYK9hpv/y9ECNCLD+8R83ke2XCTXfXo
FTiRUq8ghRYMnyYhXhmObYjvEr8yRbYvEAyQVzlKx0QFQ+xaRiGOk8L4zPDUImhzS+BQvgs7X4bg
cVgm0EictWP7+XBOH4mAfeR7QrQ/aigQn3p9qPVC9DTjvQ8oCEbPHZH7fDscne8d7gSwclazVa3a
tUXj/9vO7zwDLWAg6lrcJW2nYxbwl9a+2me7qNMBBYe6xNqIG3FTPD4+agd8hdRIM/H2vOUYYovi
nJkneY3hCrtHLeqM5RluN+A7e02QqwQ2260LXYDUI3RRpZQfssNffh0P4nDq5vU8X4mMNAXOl2Px
aNK9ztdUKXT64g6yuPWCD1PWxRTpsMmgGGFHD7G0dYGHFeBvBOyfjA7UNv0d6XUUBnJJ1Q36dsKw
+OfRw5vP9knFh52KPiYZ//+RJdggBm/eXRg/mCaf0PwafV/dLGmVcSu0VNLcPWl/RcMAvtslMUG5
GLWIfj6cwmMC8ogcT8BL+2F2PvCe9CCc6Vv78Utg1bKDezWSZPK2OVWO0foSJs+d1udb+h8ndiWT
mHc4eR98aB73wSnyMhMxg9T+lThjEHxm+VdwhSPaa9VR7c05M9r3vGHU+XBQbds9wkTh5WvAL/Sb
JtA6Wet90d6PEF7TEcjx06G3K7Qkip9vJhAEFxw4qVZYe2VqOPgiXXamw/gYNvlTNKKXaxaqV5mb
01RSUmWAWh6lJARGqOREgVCNKbp3DpMS+P6jSvVRKzjKtJlITBXnjY7cS3iyVa9D0aDDmLUVdt8L
dT/PQqaW8EpL7xtsu6RE2FUhuJvCdGOBxvrIhGD524pCnHqf1M06RHo7TMANXeTVYF28dIKnBcUV
1bUSiBfG0Wy4qcR6914feFIJqxQ3/NVD8nStCAlVHmiP3vCqmFbIIAgad7nlXaJ9KmcxtOlAjzx2
j5ZH4P9O2IZKBHIbjHQqvYyc7RW1mBoEwQijai/qD3jLOr64WZV+T62gzzbx7//iPvaMGAk3lrZ/
JzGvYdnstahdUq0l2EViInscjjGkmECzTgwoFti1uqQ9lCFRA4Q1bwEMNhzPO+Y8dKcraUJTR+jS
iFZJbEW8Vw/a5+sc2IaCJ7WiQ33vWlLlYePSOhD9UaHZz0bE4jNaXgR2D8lruLd1F+iJ+GDcZc/L
/wx6z9StkhdkYA7EC9IWRcEC1icj8BOiVumRMoCVEWkS62hCWhUCy/QcKvTdwWN0eUH3gDZ5zWnH
fbzQpQjv6yF+qcPnMEy77VOjnmAbX4psZVr9GojbwaZue6SoJaJv+/4xOMlA1JO+YKZHE+ZXj1VY
95+9z4+pDp6LNImvjZZrb5WnhdeBDo+aAWfjYI48CsIB3wy2PYfR45qZ7/uzJrJ/8Wp7WJYrc92R
TjvTEhZ/hC03LC1AM98gC2MpTbpDi8vclkNQZ0RQko5GcONC1n01bjMfjZbkK5QYFc16comnWyPu
QQLsm6BTpOQ3r9t+cEPIlH3jC2kaf0ej11/BXXFwogy4tqrh5CGBg0v3GdW1IXQDR5/4V6vGaq8w
duvPv7pJMfz9gTe8dCdNIzymom5xsgVSGq0DntJvDok3T7lHJxQ9HbtzATeKn54xdJHP53ZuZZ+v
Leo50FL/zWgsxTxbnmeG5g7JRsn85YPLXL2R2FM7LBtK22cY1g579UxgX29tspwIlY2fYFT2fY/a
k5smA4Mo1px8pJ7TgBCpzBRFYpukMh67uFacwm0RX6DgWPdbhebqs+af6aMWarzYIM1iIVKecEpr
vkcf//LxJ3Ha9X+Q6iwBlfMTACWKQQzyI+WJcp23/tEH7EuGGcq0ClmUgOtaHYCWxjUppPyLZhZ7
9Vptw3MjDk8Z46+j0bdwmHkBMWzN61TuBg0VhES+iKl5WP6KBxdF9Ynm7tiEE6+aoiBNYMPqf+Hp
qtNxaLL+nPeBLyPBVaHRzNsvsijL2QUB9OWBILLp+dIrDMSaSBX1FddDRb/9tqRBe5B1dShqSKEz
kBYs1ufp84w9uuLW7VC11fA47jbBME+QXWunL0BBDZ++GnGYboH/FynsDCudohR5JXA3Jj4cNyQ5
0Dz+b5iWm3SYIhXqzzs3+A+tojp0RJ6NLNtLaG+E6Z5A009oDuCp3aQyZcsLWD3A8TZ0ldiPI7kx
pNyfhXJZrs9q4CUBOZ22yKQuMTeGdi1Ol8BTIgA+DKIX7CDeOfQ5oujP4/i23HCJZRNeBZjZan+s
SRp7GYNcwzKeD3lW8CBVv+dp5zEzDCsLPn/Wm6wz2+Ylo/qYYfsOOyiLAyRTL6gYHOEPavLqB2Yl
RC2QyxasJ2L6LUopY+2wGYRMHekE6pJRhyBqupbZTXJ91uk6xyQtPy8EUdax7JQAxnoKqpMNjZpg
nUc7joOBiPvR9YR+ZHqk9BuDytED8AQXvqG51eCjKi69IK02UKzC+Y6NI1MKVgLcBjGD06dYrfeo
M5j7EtsY/T0z4UtcgcmJMMLjtEwYpB9CS5+TDm9Sk1Mk9RRwpqP8fU0KWEmvLuLtXb/BUviwTamC
+tcuhYtv3x6BGd37SPxPa2rxuheHBuicqavrHTrJAXBXNaDXSTnJVCwR4CihrvPiOcSpXG89PZ+/
bSVPjuGVpRHUU5FIUMuHQ2xmBZkKekIF/nCkwx50VUGmmu/0dvwtIvzNiVlZlmjXbVKHd+BmgONu
UaT6l8ZhuOCeBCzeWp8qnBytY3vE80GPWr1rIlfBnZxpY2cT9qGquSy5eiofIumgDMg0+2U6JCnm
cQUlniYK/cwC6m7B0eHiKxcg8RYZkhDZneNuwLQ0lQXSaBuPz4jDwjRtxPUqNSB/dQKAQxboR0Kt
egQ++JqSsY4d5xEjuy2hcfn0WToCs9NQThSKwdkIAZee69nwrd1M+Arzxt5SxUrBgiGiRji3wTSe
VTaZx4t8TX5/LSuwPF8elIU9ZTp/ZBNXoBhCImAMQmO+IIzi3jYF0OcOEwYiUBMvznMuh5y5Vo5y
HHvVufoOFnh3ODfA2/9ZusiXHPpZzSKMHkcvY9tfnHvvik/LB18LYFfNNMl+uu1GyvbvMTGVtxyN
9yGqIEZ5PbXfcFf8Bwvj9s+cMq1al6BFUqtsXt5FtfeLTh3wo0uxPd6xwrHbIDNj/qUfAJbahUxH
fZcd3WI/u2hzs0NkWB4OraX/nR9yK1kWp/37etcLIctUZME2lI+7GECwWjEy6c6XicMcD8ugPa3F
7PyvcmfSGhWvrS4bMOCcOvpOWnmoEQrTTYjWhgYFZ/yJT93kmM+B1dvlIafpF/Z31Uk6jX7G21gW
ho8Hrnf4tbCuzZKjhdjet9GBk+7Snp1E9sZ05VH66AjTWBAEQ9iK0eZFbDjtp6YTQAMW2yA9gtUm
l2bFGsJKru6hCRsfkmkIokdRgjdSyaRxmHZQFK6Bjt7BFj6nyDnUIO5lxCduSVq2Z6U7u9mNhO9t
48VF2+v2RC/u9Ogv1Qkmjwu7eKWcQcoqlq4Qgrq3V9chlUlGpKqgzmNK5BqYQVrEop1eZHBHE++T
915i9Hjs1/JtdabraoaWo6SaJATj1pUNlnsXyAt1nr4SeDBEJa9eOO8IqT7pBw3z1HOYTGcXrRQv
+y/TwAs+SFLesVV230OOhkvE50FgHAiODSPCVGupejVa2ousq56Z8QvclW2/OIAZrVbvvioYXFoi
FM98NL34YKzC+34XpXi+pZX5PaMhzoJS4DJWXC5TcBgiTH+j+CMzna1sjICd+Az3bTbvJ5N/3TOl
XV+lNAFwU92YXc6T5ZYomjqhQEFSUFp96pcD0zpvPBCmJzp9l+ShjDY+SICoYYPOkjLiQtMaL1uy
zJlkGCNTe/ExLpK+kOmBWlBq3L4tpSkKUR/tFADnbaNHoKiJaH6FGGHK+vA1WEqJezjwxtvAOwtG
jLeMAdNwrwsfC8mkdbhC8tXHHtkaGg71grVtJ7mjRZfMlaYdm2tlvJU5iZ1LIc43GiI7tJ0PIBbx
C9JVheAl3D2x9k12040sHi6CHjk77fB8dZ3azvMgSwXxhfabZZMf2weC2racIDoozWowmYecA3V5
SNnHMCGARJhCJq32TLFb4P//2VhwRjAr+lPIALfgD74KrO5UOIGMikS7RSMutTZK8eNYB3yT6CXR
ZbVRICz/o8YlVuR7os9iQmfK41KTOgHpwwcnCrNY+FoXHEzidp2sIyoP+eE6ZklS5h6fLJ/u4aRV
dhYqEgTxB4g7ItmP0k5lb1WwCjV+REVIpwzVKB0ur++8Hx0AmDTMd5mEmv7QDDCYKJv699Bk6QNF
Mk2pr8WWOHtL29g7cDrYZrT7xbMmnDtsp52DlhGKPWG4XVznCbZK1gVvirSXQ47j/NVocHujgjOy
YlCxzlozM7K2sAVU4YODTDnL9yTKBf5/Fj4+C1aZp7Wtbjxlj6RNnpSt8chHsdlpd+QHLtR0r6i4
UyOz7Z6/RwqazKsvyY2qOX+Jsv1r/uWOJQspvUX87cT1SdAFJyTDU7YsEA5WTAzwOkm/UdTnih50
sGczG5FEzUvklGxUGGivrxSB8i0YJoJCtCt/9Dev9oVVtry43OFJXeMTlRxJpEqWvdzE/zf3g+bb
DuY3SZZ0I9EFKxxyrrpDM/RlIzvK7aiITxcv0OgTJzoxmn6zH4dd4mgw0KuuhZUV+Q2+fBAInQSU
D0F5Lp080R6AFs0AABEfdPLQ5uZs5foXY9WlVbEsjxNleS5XSPFXyVLV4iSA4solt+ONbPDrZusH
FKh4ffEc1OP1V0IG7KTn6Ze2wuDsq/2EHGKFyWdEGSvAbn1Yu6kcseJPPoJQrt+srRKlKx+uGJfh
j4lw6OWzYgl4DOC6AUuPRZs1kzIGIzQ6sqkh/OuW92ibV8BDHIvRsmy+N0Lc90b041NwJv8HE6N2
96NbKbNRfWRYQ7XN1VWwmKurCTTECVNFQFD5ANQXs95otJIcyLTtaRuSGcO+iY6L+2Rsxzo4Ez+w
WnjurTN8Rabo211MTdDPvYcuibwH2qGSydw/g0LTqZyFHaHpnqx2SO2/T6TPspZPtTKQC2kxkSr4
B/VTDZJSNi9RuxMnTOAMG31m2lYTAQZ7H0B8D+AO3YVEy63T+r5MDVyrEhWb6fGGCacxB5g+B+T0
ytI5DmTH02waDVnqwzqNfg+PzYlWnL0DoiiYDNIxNC3p7UV45bWSWnW7tW9srGEzNxEel33Vrg/9
8Qx9IkLW8kttLEP4tff9yOh31ee+HKW7bnMrXump9gyt5TdHboJevB2JqNpaLQEHSf3L33xok+1s
G1n10q8LEV/I9GeKKl1b8NF1cqUMWr0JUUK95F6Nva7eOq4sZ7LU81MSsIlG0m+o+2wyfFIUvhID
q2vuvsMTRw072Q180rAspwiJJkL/tKrKsUm9gYngHzRWUW/wUbtN2oZiMgE37PG2TbTCm7ygfowy
Be6SryGKdwU/WC3J5prza9EwyEbY4RvvMByuTZKY6fK/IBalL6uuclyABClu40KsWvOEEGV1TuYG
pQWgAR1j5N72FhBUigKxToKWlCHP1MsBeYcm/PWNXaU99W09Ve1L0At2wKc2E/3/yMbIj7PyT8r1
xcOnnjbnA+PLODp8dksG47eiVKoSHk02ZGHEUQXjZDiaYayEkruIb/+q1i5ig+fhboXqFsqfVQ2e
I2fqc7dPgrqbRgn5i64z43s6C1zOUydctIhvYK8G9JlyOIws14IxCnaRvO+H6UJbcikPlymSKx9A
tfmU4YHdc9DbyvqHlIuDU1/364/pxQoqUcWl1s8+W5L/zMh2ly6ghDu8WmNpG9pdBUP5XE6PLHzf
uQeh6nGtY2gDxulUdMvCKil7Rb2iG6ROJbLaAfJvE45VJRmxCo3HlfxsyMjhRc19rFVfRhBOXa0c
MRRA0xfrqR657Bxl/CP5FVzYyxaWdC3q/bPsnk3clWRhwYWg6c0a8Htja2a9JBtwoc6SO/vGGK2k
IG+YGaCTPUzCgywgBv//UqTjq3mlFQyFIFq96TtDth8n1EapkZnewdoY2N4LOYx3m2WX+Q4yAoh4
4WYNNNfs9tsCqFXnunii1TAUg1/Ks4nyso+61F9e34FdEx5AH8a836JJ4nghWxsqPUgPDQflUOmd
D8F+v219+bYlt15udio1168LZ0K+ps+VXkNvnVvkiJSXA6lWF7OsesPucIz7Ra+de/2DTtDfQB/B
EFENnlWBiuTr4Cxro/t5QE+Nm7P2PS3+vBsJdfRkRvX1g28VSviIBf1h8ZChzidVUl3QDtNIsI6m
x9R+gHQ0L2ceT+SzMg6qGPFVVZvwWFkfuhc69sr6wmjS1vfme0sljrKoDBHM6sNHe5W49qwuJT0F
/797quWERVtmaMdQOorhUXalrEjuSneWEGIW6JBjDR1CNe24Kvd5dpOa3LmSLHYo/iTg7b3ScqMa
UKwqMPhbCdQ1MDkRsKyIPQa8mbl6ZwTacSRFvoW1M4qJNln1PqRT0Bo2uIeMwqzAJ8UBnDmM2syG
ycmkcRbSa6TE3jh0b3Wik9ImEIcIlpvOTJ4Uc/XeaBiDJeoozzj9BF4k+rXgQSDWW9bQFyrCI5/n
T7Vq9PfJA2pGpI9478f1kZyTfwSgYdtNqKEdSDBkCXpPQV37z3UfczccIFfKfTiRqlZPrmoRBUSZ
2j+e7pYhd3vSNHz+1cgmhkutGg9oUSUYHHYlkTZ299lbf1tK5BKHagm9aKnnIg7Xr3/96iEaGJvX
X7zI/1T96tJq/x3go01jsvnKD7pcymV1HRAe4D03kAXBkZrcHe+ShFhUjgqxCaVt+iZ2rHGQgIa1
G3Exd7GZUfqHFHOMsAPAmg2LvjO6PwZYqUi9reYE1B6/byI4G0amgpWQqAEN/ZDuhD31PPA5nqar
be1TvuhmPyTYmPtTcdkoTNjPcJw82vD2aQt3kHMNFVWc39CucsCA6NjwBxD+ja2t6Oz/ZCHMoJIR
VqxUAc7SQfbPI8v3lP/YrqxpV2AScO6fxov0nwJwZMMuu3GpfSaCcYUALPiclWR9y/0+GvQ45FPQ
W70e9QXlBjwLvOMcH+ZPQZxmrpoPkN3u4UD7djUN/LWdUwzkDFe+3yW+jnyxnQfl3Gm2ehBJrEqF
Piboz0pN4QSYu2T2ha6RsnaM4cMyu77dgq8SZA2UwWkP8qhdA5ERHj5IeOl211zqtfJXwVDP7b7Q
/t3LSXH7mGQUhFSEx4YLegdXAT69OJRaX8L6swmyMDi1vqj5bh4o0ToNX12LLRug6v1xxtLbVjYn
k9lpZD61w1V4aTOCaD+uVPycvc2P1rhdIJ+K2stDFv+iYMEYtv273NK/o7oQB2SHpFpTwje4PV2N
B3EQ9tTH7hlHxsO0MNVP+ikPIy5v9JmNAOA+MAm7SQHt2cKITH0/l5GAlAzT1iKTL2XI4LK7T8Ms
xxMhdoVPLWEu3n6UZQjoXWfRtZoCPAeOG/hf9BQxQq1FGkCWOU/vsT/n8bQfOqwhoaBm3eXg0CZD
tMSrF2PY2UAzAO17GOSTdsL9Uh+3GvX3bhk6l23ywc13sSqiuh02SYJyZQSxhqs5QQ2o3Lb9wA0+
H8goVaNoj0Gij1gQu93Z3zMgRTcJdjBbe21rwUELYr3LcaL3doEK5gRsJLwnsqnUjOC0FePJ9K4P
vtC1lg8iNQcs2VB2d6ACamw8giQiPnIbFtFQbgpj5vlp3fBU0cjUWexzKSks/HlHn2P8N9T6i3N5
huSbVMwVM0MhRXAyBw99buAw5lCTK38Pc25CckkFw8OGo/AtiRDcNtvU0XRP7mOuvCxR8zuEWwMB
fLJR1/E8Ykaq8p1u19aEht5J7qV+bZo4898LoX0nZ+b3Oa4MdLZIg4EVcZO3Ariii1fzgilmmMh9
C012Pq7x2u5KJWl7lfSWGWBUtiPiqTPejos4C/6qSfg9p2WPRCn12xN2Rkeanj4i2H2BstJ+GfVa
yDqNTVE2GJBKdizHXHYVtA6/XuvUAz7m2Dj50MszkRPGpu1M1mrvwsT6QyNB/xQpV5ZkX9wmDmBU
pnZ0TORZAWBwQx/4ZkDrVDP+rYQ5cnPk59h6FjeybfnfMlEESuEO3rlNw6BuEmE0uyuk5nV56+ZA
bRu+Eh/aVvK9IE0RBgEQMcm8BeTxn7SePv27nUgniwJ7aQXbatoylzNn8buuls7hGOG/ty4U0e1Z
G2KvlLiZj4EiNrQ7qCxMX+9tCrgYff8MOEYVPMKzxm5Tz/RFklfHbOYLbS9CHrrfcjYKPAocHsLQ
4LenIUwNRvsRJiUp5eIruCFKan7aaLyi2OS8f3YExAAFwLQehg+Ka7xgmLAlGGA7g0V/QLvynTR8
v2qZTt7A2diozkZPFBgvnjFnxVrLjZhEfgOv9n+NrYxMpMTr0DiEO2R0DRIfi6tmrJc3qjYsLA0Z
JZn3c3ZVdroouA/QeTIQUXgS6bqzNKEw31IgWEndhRtd1H8/FBIsumNcwdsxAxe8a/z7i6F4EelF
r1sKbo8sH/i/berLgXLpVZluhej97G/161vyjEPAT4VTXJ8vVfijcOZdxX14hHxIlvPbxBGzmmxB
Rucb/0tsJL6fHy1WLrIYdbQtJBQk1UJToEvS00ojaUBZ9nFyLKhuWC1+vt71RhLkySqObWx0yoRT
WxcWTfI+ijnFEZnKd/q7TB/6yo5OoAPzv3j67GIoGndIRHeJ4gEkp/hhbyXPh+pqCZUleD4XNgLP
V0tMuvj/Z5oawjkMLbgboHCz+HAL7NpdbHCKPAhhkbYCm0TDMpC0MTy7gAUOFKBxenidhThyaPvY
jdU7uvl2GlQVZdJwwVasTRDmOFiT2bFokAkYpBUScJfh/EVxVIhJgdXkepFdUv0GqoqeyBXRR77h
Dc1LANA3lGmzWnvo3wzsp7qJH3iATakXJJmzFrgvJOmtRkuTjv1O9oMzdLNLTGjhkI+47z4vkOOl
rH48h4dMPxws4c8EprUucahPwhVvd/M8nbZ28LRrTjLsCsrA7iJk3KTzg2NjksxC+3g7GTSO4j1k
gllt3Pctr6G+98YOaJ9ATAw8Ru/hf0TL3Z6hUjmyb16lZX2wuWgmA6BpoNf+TnmsqWWyEdJrlTAQ
3gYPioWzUVyNIVyXOJPaN8bRyIcSsX8BL3TejfxNAOYKyx3o2h5S6jNrdrzR8JGJJJzwlB/aJL1z
Yi/GNOX8MQN0PxGReTZYDp0boMvGxeEUdazhosgoh2WHrWXgOTcMLbaV8VUGFYLmyfPyVN09b5VR
K9rwgdkSM7aZp2vnT54Ei/3p0oErUBbmpTbXlLHx8CC/WT5zZklOqPw9UHbExJCPL13LCXoygLrz
vsfY787F1+F5Zl0l5Vve3FYmdJziO7zDNhCEsATEY5wqmxkvhp+rMfhvjj+An0x1u5d5JsOWi7BY
LKtKECe5qmOASC3WeHOcBz4pIlfhUC44CQIj5m9cKl/MCnDkp8fQccOkPAnyTQS8X1a6ixqMaEs0
0ENGmEO6KFvrHZKDh9NL6uJnHKN8gHYu5NaaFmwxlKkQfrPv0l1dAPzIBcArLzJCOfcyC1gKFIv9
tXHL6rpFXa2PEbaXG1tI0gVRFf9qkg7q2kyrgGYBTNvC7FFzuR2MHvFpJ8Vf7Y3c0t2BfWF+Sx9v
57nOtXdrVgjmgyiUBG8p/RNGRArE7lPtKGCarGF4lSz2KvfKNWVC+nkpjibyDQpn20wPha9Yriom
itwUsGBgBflrqWBY73r4BjHqQdZtQu+CH0X6Eu0ZiX2/OfII54mekfmOLvUNR/d/dk2JKm1RPbjN
OM3H6S8FhnYd5u+aNSRdiwoWo8O2u5w375naffOJ+iEzoTL3V/nIOxFJ5qcaOGBs/8fCG1DnaNu5
YsibQiestB4neXWIgK6Mzm3ib4OXWuBjKBvIaeKx2x41DQCWXuvqsFnEGptsvzrBDs8ME3mZ8UU2
gSbKVfLBmoOdw1TNVxq+z2p9sOLY3MKP28UW/uCeYbofKTJ+sgYhnPeyPn5cWGcJXyNMSCXiWqDb
6Rc1fpK0RJwCXc1Mq++nJEeQh5LyrDHWHZaYod01pjETqiHjfEWHXq1KRSTe6U1/8xd3uZVGBvEk
MrEvQVEDBmzuOlsc4UxP1Mzz0EAQ1RpbWHKdAsbaCiYshP7UW7dh71Hxp+DIzPeeQbb7a+vaaHnX
JHSVIDr5iR/ppNdzbXgUsHU+wnngxo3wggicquTKtfArwpegGpRclTNkQHGqFUp+OYDDryYUJe1Z
ds6jxS9k/TZZwTGSXG5JD4i+ElrQ/gMAk1Wf+kNDvZbvKb7trP3uUtPWHGqrzG38zT8R1SADLSKA
nQcqlZcab6UncbUUG7GsU10Y4+KuHSGfnGfcdhT4N59jIQEuMTi337lEWt0sh6xwO58CyBiWnF3G
0WPDx3UyAKd5R9NfEMSAMSxZVl9YQIhE6M+0gGEVxIXAxLYH/JBy8qBDClZIsFXlgdbMKLw4/quF
LDSD+U+eIkX8XRLCfzBqyIV8t4/qOGpzMat7CgND3vQDbraVmcP3wJ1g9RY5MNZ88zwnJe8tlsq8
btfz7WiZAcP3MsAR8F7E7BfPocAwE5w5LKAQTWZ4dPTrwl0w2IR9XziwbJoYVX6K37PqQd1fLlrm
F0ht8bcjR0CHixrCxiq8IKz6KPuH/2l64qg/NzWAPxW53PKBmI7/fTnx+PrYErRHCRVexLOGqb0S
+4SwhyEyHrUCmzmtUpzi37FM+q4b72n1dSAK7vsJKy4/wdDRanBsVvOCqe3ZxZ0u1xuJD6qeuvSe
/+DBnXYDx0ZnhLljtSYtHb+4IO3c2iVfdX5K+2aNwlz+wab6RQf9sxJzRoo8zVkEvxDA9nUYRdsm
o5STh0b4fjYNZRrURemXlW/Ajzfys87XX4R8MEPZI1xEleDXngmtz4SFpN/d8YWlgZrahX6EY/OC
inW+pgYjEB5ufamhLodtccWOJM+pdLmOfnS2MtPbjDYTvJpZBOsNb9u4wTDEEomAIagwF/Jnt7i+
Dt+SF0qG0YIIv5MeXXDP5vOwbhclcb/1ClP+ga4u+fQYDzPJzk84PjgS14yKCcum1ytwy4JT4gRe
pHJl9L+Hq1H+OeJfgJCbC5/KhhzoE27j+ponqluK6XbpuS0nAgdNj8EW/MtJG3p2hX/y32GpysHl
T+B5ZkOrulvILrGfHh8MgPKAD4RZABFSXqSj3xTw9JuJIxnFP3571wF2zcreS/P1HwxE1YajZl64
v1O7+1rHBONQYzWXpY7SjFBm3J7Z/Gjj+hc0OMkMiTE5qmuc8x+lnOnuoQY8dY01iidADmjnByf1
z/wwJ2jEREtQZIpkhB2ghnBzsoJHNBy8OKQIxm2lWysYECIQ+6OJoimI9/lhffhkJKAQIQoBJH5f
d/mH+jBwQltc0h/9ug/o8tbfA5ictOdlpgnDbP6B1xoPrm4MRHuRjti6VxrPANM8V7czcN9u1FN7
+4FjXa7kmfWxy/sNe7zHysMwp9B/2gw0OSF8t1CgVGQXnO8vAwvJ9RfPI9d0OF8cBHe3nGWClgQP
QeQitOMODBtx01WZbzqI8k+x/LQCL6FU8DiFFhvU4NlevMc1ICtsKP6hL83IpHOW64tChnP3N8lx
I8+30hhd87VLY1YAvuaDB+GFfLc8Cwm5aM5ZOid2Kx66sLCPstOmfWn6NFJIykyTVDku7cBMxuWC
6NKpotObfsrc497y5ORUKqFWD2QHYsmWv08IqB6T4nb7sy/kNWcP7z8xwi2exZuA6+LV6Gq5YVhM
84sBNqalj8OiRcKMQbe5CtzkKQVVx/F89rTpJDeiE3p24LX12f/lRkUjox6BM5kN0GBOLf5zMk0n
ohRIutox7idN4jSy6k7HRB3GDl0It6ir64sAXEO3BJobfxCsAShT0Z+fXun0g1M5bJ+qMYXqOENq
vj9oRX1P5N7p7gaBqYVC1I0y8E4/WJx12F6+y5F66+Easr+JlGh0WtPy75HQEmUzs393XLJHvKY0
wkHarwIi2l5x7RcqOGQE6pnqbtEtd2CDCYm8+Z66xqri2hnvWmicdO+RaC2St9frWFVie9WVwAte
YPP0vO8lKdioty4fcerd5LZjfP396fzqaARlEqUeuJyR78Bn52fXD1IKrCYlQsjUqwvu1MXNZiNk
e9KNz3IpyVPmAVPJkNGnUSOrlcTpTekrqXw579jbjGjQnYrL+Drqek77lsVIVlYJmXX1EoyI0Rpd
fMegOUbNvHiITWQ/g2bMjnzZT46Zwnwdu7v93M764S66x7FIS8FCmQ5mEDMCILgj3f7GYqOfFX0T
8vamT6jOEPJ0pxgTM47aQWNHyqM7mDiPXsGuibUUgx5zeQ3eMSatwZ4g8MkrABuNGiYKTnUPi/7/
QPhaa0TV1t0F2smzB92ibGt+3PncXkobWVvjAjM6J18uIYmVTDVwlniYWSM0WSVLqHzrlt2XU2LO
PbAHT3rs1vlSaYJuGVxKxU64oGX9O4CR1irSwHMFnekftehL+02DHo5q2Zncx6srWCM1mALOY37w
52eIL8IuMkfw33ht0tf12kz1UhLSAOjoTdykytok1RC5vC8NEEr539sAXWd+fsdZCk1/eYv9RnWI
W7q6iYw6vbt1IkfkD+TWX6g999H8ygNiOt1ZVsWlMre1l5OHN76xXxkvMdylV8rHj+LuchBVl2NP
Rs5dnvVrLJfIgZhUPx4dfPEJngwmz0XTO5D4Mo0JUUm1m+76dKvNk3SQUpSqj069D0h2BB1iC3G/
UkfS91krCDWJGdInDsfjuMJNM3ge2gkey9dfMv77pnmChZQw42csQkiiSuocgJ8VeImmokJLLEHj
fIEhVr/1CyzeKQ7Cl+Hpt5PG87Um+35MRj0ZlRFDgh/0lCg72zaONv+WUod9QvIduWlwEepufRL1
fmicn0Hvt6hCaqOR2xvRP3hN3STBYJG0cjOKNDC4PXiinqywke58YKHU2STLb7KdEXao7NLqTJI5
JVQs0oAZxpOXjoNLB+rgkVf9WF8FOiM2ELzWbFc6S7XDKuQk5wK9/fY3/+uTHjnCedJd/yonEM0m
Uggd/osGd7yFxxPOH7lLvC75KywdoMo1FpfbyivDZPLGTacd4gVr28r+meg05EEXVoYwdolVoDzg
STRqFcNSZurq97n8fpQkAv3UHstnXRmNgoWyPLkieHuzM4mdltP6jeiQOAt5a8PV62FjlwDnrdRL
dRjtiTrA3k7NHmQzwTS5k6oCCiXGoxg23g43r88XZjQe7s0HqeUbqCasUg6fS5Ty0dfUPgxhdm0d
29FScLZTWKKIqHD869qI7pLG80uPdokZxWn4LyfMU9nqF9FtwPQUwPq44e0V+3Ee8ww7WsBWADpS
fFAPgnbppp8/91tYtneWitcjS+7PRj2BMOcDsMJdj3mk7YLZUntOsHTDTFR0/fmua2qupiUUoKjx
ZyaeK7lGjNdgCUjc7uocwe1DbMXzOW3B1IdzwvoJrELoprgY4k0S6rC/iPXLUW0APde1MUgYSAmt
0NAg9HcTF7LaUW7Foe/Ca9DfSKNaDv8sIcuVrGd/7IxSw8SuLJEm1amQTFkOPvqJrX9aLvb5JI57
vroYU29IJpMczNZLqc/kECy3m6jWPppKgv4JTHFZ//3lqt2ShO5bp1yLwdT8mKmTGb/flpOeG8tr
lX6LoIqk/74OC/KdBW1wLd32Ci2bIzB0M2sKVyUrvXFyZ4k/qi8lHwHn6ZM+jrqE3hgJ8+aZYHzu
s3dq/SX1jYLz6iwX0yQvXTGYAeooOoQQGlylY+X4GLz7l6Iyc7Lp/XdRCaaPpZM36RYZ7ZaWn79q
xUF2M35c+9sdUP34geg40iB2akaNNhnlDsTGpQuN5bDUfKJx2diCFLvaPUykFSVRZWe1GJWC95jU
InNkSrK9aqUN9Kedu0OVYP3vc8RAVFXptO6csOd/le2xe4/LD3lacwqe8gnfFIMQMFFcl3Eii9ZD
5fOPutNKGZx/nVAVSRPgtmJDx4sVOLDKStOtONU9UFMiBJTCNZe6FfWPP4aIKIY9BEf5grzsq/Bq
2+SYIjYgt4/oRwvX1W2lVRE2ERYTwVRhIhHMKE05OmB3tUNIcXseBVbXxoiCzRplDZYLY56Q3IoQ
tgPk/le2f9GuKlDLXVNxS0Q92NuUwT+2f3NX1aVT8bmBVLjkyK9eGl5V/gcYAnidLQ0JI953C5AF
lo4qfXv6ppJyzCSfpNaaVeB18aq7uvFxW4jVMqQm11HNKPg9vGc57lI2O7A60UHYetzBDDFDwUjB
GNbLEkn8PS9TWCi5NLXyMToyjLW9Kq6/I4DseFYT0NdCZUpGckaEJ++HqniXaWppUUtf6x/Dax35
CD+l1R/Tz6X5WRwc9xjzn8ZRxq+PjJDvO5Mpw03o3z7HCDwjXLOHZS3CmXipFrq7o2Y+0yWUUvSM
HXifMUBoZChlrJS/MYCkUQns5rB2x718hRoClY6bJqc0BPKdRDgymv49RTmx7Jiz9zx1mvB6Opc8
Y1bOv5VkcCGAPk8BzDeLeCHDlz/APjS8zgJ++EXt1FdMRTbvV4ZlaNWbTW7Q3yMxCQSFGcF1Ln5u
MfgJ9W2zeCIv445yLqYlKiq2td7riox9q3uNlp/TaE75PGzI221hJlLFdzmKs/9+HcUlt2lul9To
gjY0ie7+AcHrn/8YYJI6oLGDN8DCk/PjKU7dNDaCfK6bAU+KtLurMPdJwaUVkKzRWULSHIC0cwC4
oh1XRZd+RwHLrpBOQR4diCi5yGxGtd5ssnzJ0ExFbxh6md6WisVprDtp1snAAuTw6N67d20NOgtG
nGESNi/2nLMcsvDeD9NxQN/vtDxJ6zKGOGIMRiK1hcsQT1rQ22IrRpA11KCBiHQzXUdqtICj8XZQ
udr2pbsKc7Q7qBjWqMbu7aCb2Cfy+VJy3cOSuPAw8GpL7RQI6DlLfOYPSCpkQ+0l0+3w2T065c4U
kctyN5GprHodv/eTWdR5wOznOXKcd/aMrt9b0hbsBTVwq3tL+52OlUgwBoY019riyK13nocGvAL6
1C9D7Z9QMEX6jJrNj6+Yrg+dKMVSVjdiTXUEz8FFpJpYbTEEPfslNf37D1tvs4AEVDOkBDRImNCv
4flDLEsE9GOCAjlFD5me/7VfwNaY5ZZa3XQLqmtkDnRLsKE56CoJD5xNELxXu7tRNOcCnRY6EU0O
2R6tYWC5ICi92ZXz5B+Tq25Vmfy3QNvFP9Zdb7Te7nSpaZacFBi1VsMH4TarBidla/b7VtoeSoOU
4qnkg4yXHnvOdk0KkuhnYofEDAJykrqHXLzv1wegB5OMJY3DIED0qcbgbqEbVcGXniWTLmR7wfLX
mZX+Y1knbwb/7Nj7ND4go2V+I1BH3oWiJRk6FINZI8KDuel5weS3hr6/yg62YMGLFp0gL8uz8yL2
CxLYWvmO8jnSkcljuWl4KVK9oVrdNF8sLVcJNC1aeh7mAgG4VP13GByFL3jolFCqnXFMNvUrn9GB
sf8/18MYj9oKS0QoYp0WBckTV6ZEf8PBDqD4DgmFzSTj0Ba+3X5huXEc4b/XBgAH6FUnIPBfJN0t
/DnOSnd8bUWUdS5kUsUMlg8pTnWY+27hUPP6tghp+34IthYj7o6fT0RZAW6ncxa+oorSX9OQuFlt
80u1/DfJCgjRSWPtmlFb7oITePqYtS0OjPX0M2RHyWFCndTBaqneNX+J4gTDMZQMyc0++EvF82jS
jKsKTedaZeV8gPFGTYqfvisiNXEReNN+89WSRSnkb4zK33mrkgdA555zg+JDnkPO5g3X3F7348Ff
0ibyZwMj/J62jbQSlvvxYKMNV88dY+v2ETXpVpbDmPhqBDgRuZ1lVGt/sm62JgNGa+KIehMW4206
CT3qDHZoiM2MC+5pNAv9XIyQM5VUtpnRwhtzGI7xmUZLrYnCtvctAqPL6S3xwsjKT5FVqMzQC9aR
Qt42NT4CCfQWoywzGWlecmU6GCzVWYnGbixtaddNu0E0qMzzZ3CKs3+QhjNZ71iEZRy9mfMSFCrR
/nRch1wspmLxbHhHPUO/kTh1GDOMjetpUgpkPi0eL17n9SfRIkvructTtY+oCh3piWQ2MFvDorLj
Lsouhu5dL5PtY+VfEyq2//S+DVKVQiE5o9q2qj61PqWqti2qg2qYBGedIyGL/7lfZSpQw9G9FBv2
8GJwxCNnUDnzYTUPU3DTdpxsJFP2sJJwYkXizOxxiLujp8GvIjZ80YEeSy/6g7ooivvPRkmmwT+X
sm9/cUsaGqDFuafpSOMIl8WCi557yN6mPL2PEc2m7WJHAYN8dqZEvpnmlLiIHBfKxLRSv1gbfGZJ
raUMFXsN2Iq06ITsYMsQp91bmiVb4c0Bcv/j08S3OnivYumjMbB2ZdcRz1cAAYRfhPOcd7eK+GHj
2vt0clsbRV8IK6QnCJPs25n6P9mBKyFm8/OpeadicDWBrPQaNkCfxr7ogq6zoczaDO6Pz584jIvS
XIxu81GAfJjLL7nN1hYIGOGjIcMUEztK+XiRMJ7hDh2HjLqTngfrF0Rjr7Lkfw6dj08R+sZWpDhk
iSIk5PvNtu1h9esWPl8wOhXTH0nyz2R7E8XI6gPdWly78RxH3wVOEVx+VTHdcHRPYrz4A8932DyW
XQUVFkGcIztaEzVURjwHljMKGMOOw+cdBUk4KYE3seJBvuqOeHDqnSlCTXmjWCtRNfkrpgxwwB4V
7S7dheHkrWdi0J9T8FyPcqwrB8AV5OAUpinSbmDR5ricBeey1yiW4LV2wqjLmTO8AgpGxiKazRCq
ZoofHhDkTGCaLd5E3h8cB7+oD+1igE2S09wx0pZOAvIvUzBA4n3kydSfjE+1kLHOhQ8pBowHp9A8
dZLw//7VPG0tGHXUu3CwEFwFb5w53rw9MtnOxypGo6Z0H0pC+r5Sur7X/q3rxqzp7QD7kfuUnyT3
zzkbjSsI0Xyb+bkL0hmAHoDHcr3J2Nlg/2rFlvwRpNClaT6pvXk5qhvI4xHr1pxkGPFRpbeVzqDq
yIlUgzHZgnvH3GXruIjSrOQhw+Sobku6AKf3+5iVMo1RNMZq+/lo5npFQXGLtDGc0wHQFttlE6F5
G2xE1Vma7FUqQQrTYfzmSJln27B+I81VA8Wn00tRTQISzGnVC6vdDN5ykwRjbqsOOm52pBc1qbx9
T7+I8NQ/MqwBIDwUNgHmooezNIylNK8O/Z4kVq+YN6wVqyooYFZj/mdvnY4bacwVO8P0wO4uiWPk
S7/r/QrAwZLWIW0qEY7AyXmpNM/dhKcSbJNOoyYMs+mrVMARDSxHATd4X1VAHoXoA/TQEzkwlkd8
/WZNHY2m4E3S+fkalAnKdOG+1ZY0Wkv6fnLu201XDsLlgehndihd/h73j52vyOD9yrJajjD/LZ+J
bQOUGOdAJ9XUTRk0OkG+y4CAK8JBvJo+ueHc0rl0OcZaGPNrH/+BN9qU/aRGiQZY3z5GxFMYyB0q
M5CODFk5p9Eo2AeX+OdovWpibqptswzYPy9puJncO2976kOOxBaC8d3Tz2arWHBV9+JrpsdfYHIL
ny6njskl5NDA7nBUc3XqSudPmf5eUip3zWXzku8cw5oIUUvrS0l3VyYYK5v444x2H0YbdLELEr0z
6FCYzIvzP1CbS4+WTUGapjFQuMxX7cEBSuDqgnJWhgrrDk+8ywRAYAKl8J/7T+T3WdJDrhmEgyRJ
UZ8hGpO7gEFxtECeCCygA5RCiycd7LZ/mHKZ1Fc8MT2lb1om6ov1g+D3+ifiOD3lvHcpWNo2U336
Us5TPkX9iy2+ZR1fzD8d0yO0Oc2ufiZtrVO5jMvdPlXE3e9pX1+O3gRexbPOscUyb0BuyBXK/+Ar
Hj2chQiNV3T3aKs4UcWQwCBagp0bbjFwJ1/1ydfx1Tqi3TV71gfWVwKDrSEwDWWB3ysDRxzKYCGo
7z+Xbmyg6iWC+W3TK5PxarVtjwLPH2LcQ3NEpjeXIXWs6lL+elad1thtumOUIwuTvutbevf8ihRn
iIscIpJA1HRFaZcFOee1hnl7znKCAdNBQJL+52HgI0FL1DG/ycLIyhIl6yFr1OCup06mDVAgcxFH
ZDPnOE3+6ntdfr41qXK4eJahIpskj0h+MjFVGh3FBNGdP2H7xeExiMIPp2rY37r+bHwlHichEPif
NlJAWp+SN9jJ9C4lrnmWCoFR3sP8aoWzZK4UfvcP3+b3CjVOj/daih/tQXC5W5qLupqEA+wgkwqz
E+fBR3cJca0H2n0B1eZQw9GpSsdCHEQsNwB7P0XSLckG8XPS6to2mmsDmQJB7UdEgmyvAzrDxIN2
X++Cv4hu442qdx2KKklrT3Gw/2J2s/0yScd0syY4YdP0we9qpxpHK0BPYW+pUUUC+bZkX9FCGbiO
1AfMEOG009KbcjlMMIGRRv2UFr38u4TtCHrdHWAWv4+33CXzjzwqMzht7EdrWBHj7diBLorvGVyW
/+V+rgsqbhv6hH6N76g4gOrJ2lgtG1QRWJm+hNHbQm+tVW6oo/UBsdGEu+3cBIQDtPt+810AEJFq
m0QlF8qCNlyfXUrZKleMwE6BQKhKHvaWXIv/4OISiFKHI2D31zHKA+tMa+LTpmujcejQsopyHHD3
+H+i5+YmQCK/nejZn/nLI461NIl5fQ9IPssXiJ1iFn2t1jmlz/keMG5TqoiOjMNQhSkr5C6/OC0a
fr4IqTdMbd+DxLK6Pj0pN0XMP2DukY+M6VqlF3R4uRvKFX/WnitvrLyUWSOCRLrYLPqwYOq9YDow
WhAyI6vGCmPzn5L11f2Xu8ki/p8K2z6nzxFst2fNyxJqJBhNUzHTbqPcubLAWQGXV/Ri290h2Uhv
zjjbRzxDcNghqQxXMxODGaDS/jcFGRMRpfmU2NCeQkRVIdRUzzMVqd/xydVGH50hLt0uGRpUkXH1
Dddot50bUgUPj2ec8KOw9R2PrNfwL2dUxCu7aetwWRnO4B8pDQzWP4eZKpdgJbNiQNuzYcp+ilio
T7DVOluvGyUl5Y0qoRZFQ6kFBVdc5w6FDOApzlL9UbU2E8xclmNuW85oHLrmoA8c3nIUOpnJqhc+
0ivcnliwY6z6/Ax/pxuxp5O0KcoM6hO/P1CATzZxz5b9XV8URkm510k+HOwrs2vrwy276KPAFyK+
kLsCXIZ2TmWdsJPMuwiuk2cVPtADLlX29c37rcDpG2OYeIAYBkxDJb3q/UugGh66x23B8I+vAaHL
kK+U6nogdKSzzUWex+iWJfPqSnfj3VLWwfn/Y04oG+tsQ0STqOHDMvpA3aMQeJXqvpnYm5QRdGPJ
CNA0RrMwyrjdvszGFxkT0AY2kz7PFLEViK7VieCh4qjgF5JXAW8beLrYPlXNv+0WD19OmgY9NQ4Q
WTBqt0B1/weVfIk3/I8GUTp7VYTTJl+Sh5ZerQ7tV3jMeMdaBnEeC3AHRQENJYZCDmGe1lIRzdPe
vdWIl8rUfCO4bRTQI3LH4rGo27CzEaWZrUJWmnoWG0VdIpeh0wTYSWziOTmit6wGJ20uOwHni7sY
6cIpC352GJb16QO0hsOyffT9M5sL7cSrrp/cv46aDV+sJhOW/G627aiC/SP9t4Ut3n5njTfwTGjO
F8QS0jHvFpWZEsvmxEpg25SxtuVZ6ELJpPa+zywTt4Q2wq3WIZlvuCxttIE25s488shgs8dtBtOm
nJVENb7uH+uvKGSNHWcpDbQL6pxhMo2MBsouqWoeAlgDJnVzZlaD36YXoZhPqHeJ0LNkdCL7Itsz
KBMZFBe7ToaUvuJXX271uqjwmT8oZv4Lucr2eh/qsdK20sNFeNLEZXJMY4PPkYHnGXalFNvJNxeD
SDnfmiUO3bbcG1E6X4hZc40F+X0gzfZKn4z8mOm2+9hUTB+xzm/KrugQPIXtQsr3uaVxNYpwmPXJ
bWGq3GD6OvfgGo3Hoz7F2C9Sw3/TUhreYDkQlJPLh0OtuRM82nc/2Tj6dz8nvBax8vVYaC7+1jcY
IXayosz7459P0gw69FPChSbwGrS+E+cHDPjsFSAuPSsWQBt/mwB8gV0NiodDpIWFAMGZ4pg0yuc8
nP7429mqxeHOEemfZxQ/uBvY1k2xA0q0MdQgeXqSL+sKQ/Zn75lwZnl/3niPFbaemv0n9G3xH/Xf
+riakhkpe+T93aEmlDHfZZFD2xA8wWpU1VADILuE4RtfVWZ2kSKah+VISTmDfKEbuadw2ozz3HwV
xNLwuM0VIWrptv3GpAPHu1Cw0NiWZP6ZQHYSBC6buNBvWHCY0vFGjTDTTbjdqNOaYaYgD7OhslUW
fMHROMkEs2porMOW/wzMQDVW1xD02EAbpawjj4bfI++ZJ40DcIHf3jBEq2+fRs8k7LZ0kuK8/PLx
O4irOaJTRPZNe2tXhbTX4wYK18BzhjA0q6o9uvEKH0/Tk9kkGmbVG8XMVtSJTql+9B7/2It0sN2n
eS2zRGkpkPxZHdd8oX8JgM/oT7sJmBtE3fqsQYV3RKT1aenluA0ohXcR4jvnQsEC7BDaveJ2WaXu
POrfMnGm8k8rIUKLHj1+++bJ6wdSr4sKtjIwGw1AVdR70oO/CAo4NJxn0TtwpT3LC2/mGGt5ilD+
ZEqcL3ZUrNOFkfvDlXCXndWMS0qdWU43mO2sCqSzm27LlAFt0IVDMnJxyxSRTfCbUTITp2s0nBfv
TLInZh8urTbd6gin0Sd7NXRmYU/vwhc5PEJq/izfnzcpI7UJvxGnQfQIPcNnw4wQG58RrFVKjKsA
rAXYxm+c3RFuUao8DGKMeggoTKHFiSQv9ThNEW6Rg7/J1E61LFJgVM7PdjK6ZKNfbFCv5Ro9dhQJ
+l4muRgo+1JFjcqE1IM09afvIdBAdHhN3gXKcrSgJQdK7L2cnL2yzXK5UjHI3nqchweAvhflhfDi
WEpVHvW7ROuTT3lF1LS+IuMxdUpzZAldkbgOrbNxuZhJMFYTdbyG3F5ze0z5iTKnO9k6GZyLfIwJ
7EX3Pttp3uyLqFbEGqkgN+NPFDNIxs268MPyIWuj0sQzceDOcsk2DPjx4LNTQjK8KarEDOJXf90R
TYDCKbOtpFOgfQDE41A4J+oQAF6gXGpE/Hrx+jHkknualLh905BO1gHpAH4ACbe2/kgLcptxS5dT
uSZxGjxWGE/191NjPfbHzoQegXPQHwMdJX9vGIs+shvXWfB9BaRJlc6IjbXn+urM+UlnKY/7k+G6
S8O1Fk6f8CthS1YKx5C0oq7tNFuzrSNb/punWnaDAKFe/hgyFah06/+L8LdbclaNARZ8kR+wvmZH
ixUldQMEsbKC8fzf/iVgBF2IPDcijUXhICmDUjRn8PKr+ZBQcNgNxONas2WPorbksUsWRjouYxTC
2VoyBTJZiuPek3qJSHXynHmOCvxarCBfxCrZO6b1c6lrXYqjWAwsEikZ1wGojOAa/aGCkAoWNtJs
2wJdEPrG1TL9olR3cUWK7oNJOo3t+62mBb7850+VSFCEzNeQN7N6mT6U2nhxoajrAuBB345wwldu
86Lh0qIW8R1S1qdZgXXimiksOW6dIfQ9Sr6ruUBVPe02GvpQwa0oLQDBpZrKpMpIO5ZUeAymrvxP
ml6EHg9MxPdWbdAAD0rMM3EOw6N2Wx/60/ctFODfH4knqrG3hOSTY7MO9MysDh6afyvjml0V9tk9
A+pAX9em1cnNy+uHlAtf1VOgc29OXi2anYsOBOfo9iasb6v3UNx3zaMV9C71GrHATU90FoPM0dL+
RrHTbqDkpUyjWMKRKx/786dbcRyng3wIhtAvOAVdG8AhEc5vtAeTmy2HWm1CYZSLsd9wPk+lutrT
VBdMLfgiL4R+rEyo/k2kKQVDXWtSMlY/EyrsXUpHcFuJ9+rl6w+rZUtdAzEc3z0ZxzGKVWr683Oi
oQp77HCCcbU6+xxA8CSeBxi3v388UsKakrKjuXhErKgM+cuE3qw3h7NBh4C8XX8UcoPmM+bYVBTO
yVbsC45YtwMqtryJ/NZCScpTFFyTXUZz+8ewsBgriRXiZRCxsqE26r7BKWyLfzMWxNjQevGefWoe
rbnF5qahWd8E9E73f274eI4RpvhPDnYtKtGFCO1kV7Q48IAhcTnMQwaqSPkmCsEteRTjzuIpxhEN
OaVCfG8KTGrkKf78xu/+/YKWaCxBoV+MKR/eJOFo7H4d9t0B8c4LrSA0KO2S7NPK3UVm4qJ56uP3
wzBxIVggIhjwWS8zkyGuabaSC2sjZPdqFKq2J5XSad4mJ8FeLPimjKLz1/IB87VgjsYdd1/3s8jU
Je6w/WkEA+E+VqndZk8r10SdW22JkAF/EJmazSacwh1CDOG3vMBQ/s61M0rz/ckDo8Bvq/w7BIlD
kV3oJvjx+i/OLV6QALzke6DaNojWia8hQmnezoSBrY8pFx/Ub61tH2SXdC0nn9kwj2VhKCxi9sMR
IIQCygMai4hI0nDSIKG0O9Yva1VU0ZNIxJoup89OdUF7hERZjSV2SD2VCKL+RZzt1h0CwP7dpI5A
O6OMtdBr1scghAvWCwKWg2WA+ToOBy9ROwCuAfZ8LCsqTLbR5C4WqFPlL80rRgUTnj/IYjhqhcQ2
r/xeumz0baAeSobG6BbdQ/cqeMrhWcUws5GAivfVweK4d+seFJW+ZlrWLCWSsF0rub14MYZ75lOI
G52SS8YAG9fMB7ULyR1x/AoyDyc+fCI9qCYXvreYyQDTBgrSkSGN5H2SAPcemBGIoEpmrU42xTsU
XJNvSIhSrQZvDnoY+l/vPtA8F8BM2+0dpGi7NMnLBRdzWCLzyaQH2B9Vx9FGbO7ZTvAC5jnn3RsE
IF3829PJwukAu1Mes71YxKhAgXczPWbBEhIpYTNn6E85PZuJrCdMVUbj8ZB1XabaBPTOD0K7p+Ex
x3ZcyUuexcOupIa85MXLOzj7jGPGkOkjt2Cu6J5iq/+CR8lK6gQPv75k863u0CkgJ5wzI31cpPrY
RPf2Vq5JcUB+oww3D7Ov4Rxk0gxsHJiNtRJGH1IvM9iP59SAN4VuVRnf/WpKfa82dyG2BWk4j+pS
9Iqu9YgsXgKIUYfSq8cS58h9nDjal5BWmiDg141UiphzC4Qr9/Ag+LxdXqpTMAAFsW5Pc3RgI+Nf
Ibo7aP/oALP6H6hYnjHHcuZXJgyT1gPsY6UW5sEaED+UTovRCT4uMkpi+sOBTQoYma5SPzmyk6q5
kYMuomIU44Km9UrW6vgdD/LJ07/d/T7h2+cMdVhYbL/SrVx/k2p8yTrFb3uFT4zojWlj2/MptxYX
j01/202pXUrwS81yrDD/+meycKL/UJvM7aUzLPBxhkYpDOEHD0+T1ZIV14lXdFU9jfgHORPVoi7g
rHWiAR13dOisn7lUBGmKQ1LECnv16wSp/rAEogXiB2601rAc8VDwnfInH25Sz16oGYyD8nUNe4jk
/qMqO7KtzD2AMJIQgVAu+8bZr9unRo5oIfv41jG/CPT4OW84Zus61HefaKVHKjjDFC6tzOThwvf3
4rJ4KqIgiFNSuyr9iRYRlLfwEeSVv6c+ihbvyTga+QsADL4CQV7PswYFJgv9pKv6hLeusg89JYyv
sGQeYySSWibalMeymBwVM9n/P5DHdO2EF9Do6wYyGAwSdI31wCYHTKsggWSCAj/4o5rntaNw5/yr
SkNLbEcSPTNI7nm2gCOcgEDF4OMECwLpiZXZ13q8sOgRf2/D6LLY0EzCJXmdfe1N6eep8vhqTt9M
EMsJ2XLewU9B39YpcIXWTxxL5JDlm1yI8JU3YfMClO1tvcLpGo7NMVa+0OBMZNnWRPWqkM/ZhaU9
3CrJTPmfJVFiBk2NdIcbgE064ESlaZwxvilJX6QtgKJlSoaWD3P6DCke9eryNG1lbXtpZeAhQKPP
8J19+EpgLh+DyiiUW+WMC28QRW9B0FJ9YNGoy99mWi5xybVVPKlwYwr4otniG3cnYOFbV5NP6lTq
fEA+qT18Vx+/PfzQdenPwkaqlL8J1ETKWEZaUKsyKSN9SyN1cjFMi7llZ34SdooNGTDSAaF5xG8R
eWFiN2gYWl8+G7d730MInjgTBxbiDsfJ130CamdZi6fQfzWJvO2AY8w4Is9be8IT26M=
`pragma protect end_protected
