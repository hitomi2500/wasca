// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rTuwIyoKtC25Eju31szuxXkuhZjmIB/eoWXhH9LbKA8X96U1mEc2UWqhc5+Tm0puMPA/J71MKEwI
QBVMrSDPkxgdAKBT0mWPY93PESbcOuqYyVcwaWNAlq1NLJ8MEqSW6ELZ1mq+N/XK//ccVZkCxBdU
iQbKAnbS/E/hGujwq1An0Hp3X7z2B46pz8ZB86YJFyrYf9GHsrWFZF7gNkZViFYFZOB1k8PWZRx+
SqO/pxq0CtdUoiG7m4rEaWafYcABzgmQynU/nYtR6PCW7RC0Ngt7RnT7lFVL4xkTjJE3Rwie9xLp
ALfbAQ+dYsDtsZlC6zWpUY9NzfvF0KO9qt4Xeg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sSJPfjFbb8F8ZO4YvAW+zPuK1Ono2gqfSjvYtR4on3l+T2crOn29Xor1OvnDOWyJA3u85Hd02+QV
sOVuMVFp/TJmL+2w5LF9QswtMNZYzgdh2r6zYxU3uuj4OmTVGr+qE9JQP5rEoijLv023rcxdKxKs
JnNK3WxBOy+a/ji/rZH7XQsUg3z6w9kGCn3zC4B5+23qho0qeOM/O1LnvSbMMH98fiDRP2j4hLqP
ruKJ0SiKIXu6Tc5BtxMqqwxsu7mXp2WeJkKHvcoiYEPhhL9NzKP070f+Xz1U8HMHVHDk0veJ4msc
6Xg6049yrs3/jPWf9umz3/L2QC4EULlp/GZezspqYlk7GGnL51nf8feL3s0g1v7RVt1bXso3LNmr
zarbM5B4aiyVbFkqd5L61Tu/aBiorV2/t9mp5dbNVtgQMvGfXmVZmyOrHjuYTHpV0of/k2WTPHUZ
KwNwp87n4H0Fs1X6s07Ez9PbYrCPSfO+Mxm+vgMf8HG+1CE8uJH4kS4a242bQ0eyPBAld0PKGqwF
/uCGiPnC797Ph3tTMStnUvsfbwnCDoI5422ETLhhuLPbBkOk52j2s66T8qQMSD4TmbN0F8ly9Wxs
yj3ALLB0PyFJ9Fs+3Jw6wejG9DpDyBlf1RWQwvC7qidqToI2to/4xWPY9pBXGCacWb29aesmSjef
OY8+FVotC7KHX0sBgO8Py3EhaFPsTtvRY0w7T88fxO5Lf1bWZaAvuiTyO5pf9Bu3pGafUJXj1T1Q
d1UKEDq+oW+jn5Slvktn93I23V5Qr1Iqh3ezvfBma/9h58W8T9U1ZuPjoF9PgeVEgoveWddnmA90
Uh4OCLSiei4r/kl4O1tccdsvFY8uFFTr2YySm/eAklPBQr6l2n+tCrq/6U9mCzZ+nsdrydiFGFHt
7Cjg7jy6VhQXL//99hh5/FvZMD/6Y9q4MbYU7VRcvFcGoXZJsUvXcr9/Q9Hxr3tzEhYM9vmTkiza
xOaCmdLeIBODz8lbW7Uvu0YTw4Zt7KcV236/DEvXrOyo2NGK9ad6YOWsensNheWV8FfJk0QKwDnY
JpjGJH0Lr8V1F/VwywJUvxazu7/hKXp5e2JqxJoP5/S3TjtNbkolCr0fhp5ZQVzDFGxchYBgdqlc
+mdqyIv1pEi28xGPUgBVBOyU0OHwwODbCkbk09Ntc/N+PaOSuGRd8VQPIQWefsPp9CSEL+lU/UJ5
ftPoT0vUQ3olQe9jzO9ofcTbTNb6I1SrslcnWZ5rPoa3tsWKtWtNOl86EZYyDYVFut+8UkFGn7hm
2oZRacC16uouMo5ZizC2dsdwpU7pOGr2ydH1ecxiJvhPRIge5/86zDYy20QM/BFZMQUyLblsfmF8
VUGS5eZzrNXsPzMQGumUxRKVb4NwRZ7ULqxZGK52gEnsVGPnKfTjmDDcIOPrr1kUQICIug8weRM2
Rgut2tLhgCjNBnuZaJtsMw2/uHdDdfYpwIWJrBKg/DHfF/MmVQyM7Ebzx5H0ZnWyY9NfTHDOJNZg
EGgGU4+vHhRH2Us7E67YXp3iRIoZNdBoeL5CWVMAQO7ugmhWcP5vXjO9UHtFphXliezeJBlJ8764
fHHw1txlehIJfjDCAIeMhUz3cU4VLQPIMWEXLavOJyzbZzsZDkdwuf02cwwudwSDhHIDZZdEkhxy
zWaOasL/bTA6JMHX7F+YnvlDlCblBFFW9VBrJR/n3UoGqLGd4Kv1JyJpsexMsWkqJjISauymYZif
p6YkYPNO9c7zeD2RS1MIPXcrF/FX9akH+DsOdrSQVk7JjszAG3/TWzHBK5nsXgbjpM6MCd/peaTF
uEfJbvYinyEYk3ivAgl8u8t9PVY8+057UDijFMoNGyTfZjecUY3+plbtcz4E1U8SHgv2ktESpYmq
uc2WSTbXJ/7kR1HT6GFk4QhO/UO8b30NpRzkl14oQsVoAHln4v0Pzumkovp+wjYhoHU9ClraIjYv
oAcJXXMzE5W1VEb9BDXeiP4UyotPktd3yZM8OBe3y8gmW4sF75NnkFXCEq6iN7qCSBHV0Xefeq24
d+JU6E4d7Cba9wjqWBus2Z5rTE3RXukLfqrjMSZi76iyAlwYyn/ecSh2L8xvF9YxYMgzhHa6lO64
eWADbVpOOQcOg1QiozXaOMkyzsKqul/VdLM8sbFGjgYuzfjK+IIx+ubMYC4LU5fBMew72fd4flqu
sq49Us4QAcJFLlQPAtHetWtPYbi7oE7gxVSRjbOvl8gQ742bD1weJFenr6VDpgujAZylan3spDfS
1K4U1YjiWVoEmMcH6ygQnQdM7wE3vt8nRssLqSpof8Y5X6JTKWTHDKtMEfqKAiWhlSVtG5FZgCWQ
mMAapMlAtMvfWbchH2DyCQXysbZIuYQQEJFbOBRAxFq02195Kl1RYz+h9AEcQdSytq7FIFNrsPd5
hN+qU2V1iJ7sByKKqKOUQu8hS2vQZIyVQgqZBOr9drPZQUSN9I/eqUaRKnTi3Swmnm39gxhmzKAR
SO0IpWo+EjmrkCZhLZi0amhVklPQQyBaxU6MxTmF5mL0oayerz7UlMZLnfAc4BnDLRIQ0JRZm29v
fIdQpz7kSErGnAF0EqFru09GZGwo4S45lfgpKymVCNS0x6Az46D/c9aVu5rfem5bE6G9qYDaRfVw
VPKC7pG5YB3UYnpmHfoi1t4IOSKEFSxNhBawXTWbKrEemLtl40bG3j5wb7P0Rpwv1S+fxfye+aBr
Yv2a1TRHUsMzPr+7pFx9vzv59r+Al2iYnsfZlkrrkYHr8nMT6klOweC8yJLCdJrnfQfXHidJbtnY
kNGwezY1tyS4JIQaTPC+TvI7XY2qtOjaQJCe0OtrVwAeoxZG+n3XIkQe2yMcdF8OGba6UabsMkaX
XXYq9YrciubrxcSV/7+J41d0MDTLtw6WkghpaS6gdY3osrc7kSqzfsLq845VJG2nlemJqsj98j44
P2NbMZJcinF6z+rkxeQ6Y65dWeYBerPkMxHT7Hcw35sMAHH+Prj29JWegT6X/NKBP12QnzPpY0jj
uuk2U0xpxUt9CFe7fF7e+CuDRZafVywT0msA93dDAsIp5Hl9G+WAB7KAoazp0qxH7b5OA3xNQnSd
sFdIt3VLyYl+y6+Tbf0dgH6M9w2VHkCmPGTFD9ZOugLsLS4q7uCe36AIbYCVZcx9CmhHA4r+oxaM
f8jzo37Vust8DKGYFByV0qQS8DmfoVU8d6Aro7QK6ooYbFd1PWbfYufssIWx6iFncLfAGcwOy4Mm
Roh/nAdOi9PQmJs5KE4vJvn14gm4tG5rqjrgGTBpmK+MXUVmM+ME2pzmmAHCZZ/Bevbpq3finpg6
50tx4j8pg3wyFuGZjoKBuZj0ec7RXJjT2pRBDYY73509JBtonHS7HN1+YrOba1OXNPxn9fd9HbIU
Jy2xl/wfYULPqeAtInzGf/FzYEaMSrWgxEo3WkNc81I3S3tWk4at+ROIcQkD1TgyL0CejTJeLlUf
3H3nB/NNbWbvR4InUk5UqZfBpzk/tE8G4x65+5+NmO4jDt2oaNSbHRx7f7Up+0bCLDX4kBqrCJXH
VvSQ4yoFRb7YvP0s64ZTuops2GXVjH1C6ukHCPSrlzP7eZLONkzqki5yRydf/U43Mq0euRHEKrHA
cGDQD4nApwNwHVppDQY3+zyi39IWKXMmPTa9ecsOrbrqQPwb/txst7J9VhtNeycTOsmkuvmT2MOD
/jHMZZUkN21BB6pVU3048Hu+K0osmjaGqjonXBauU2eykcoECbZHkB4DZZJhHpYf0ofVd4XNHsPx
rc98xeqfhmxSqdA/8/hCNhunZC77Iq6srnI5U1FoDH7Xjy9NhqjOJzwfPGHH3tr2ZeM5tl/VX2E/
Q9B4LXKXftgaoOW8tzxkKmNewSgpVGA/x31ZHPL8wM++JdlhdHWyXCQ/eTzZjmbO8wdUkbCDtoO4
n9cejVGg3EaKwUgbVJJO/QYvNF2BQTIQ/BojLM3ikNVsseyne2ZYFlB/UnwOi28ai9q950HARNTw
Nr5eqc7DaHwL0mrkGBirArob8fcLNdYJQDjlA+XE9GmwQ2nZ/madYYgvEv17PCGwj7lshl+l0gRN
q/2sKfb22isK/fA2m2jDZEy+aRS1DRiU3UrEdCcVj/4ccTitxxEIvspY1pfst0ny/lxTWfMy2TZp
br4HmEvBl+haNkIPHExwuf+h++rmXZ8NDL8yg0adpybwIKilKf7YnqzLXFMLnxUFsyi3Bu6zwarE
W9j0mkf+5LomBIipCiQoZORqLn3v34etll5M38rVI7oiWFAB+GPVTkwKtBj6ZxMubcArNmPjdJ6M
sS2z3UFAhbDrzbrpzWVWvg2o/2GvMCrV78XW4/P9XpM5RTXeF/6o2Yk/aJenhkmQcQm0Iisqq6i+
rcN5oevM5ZtSJGbQMjRe7t0Re4AQdNZYVJOHWQTdSayLEk2xHrpw54L+O1D+M6hnEmgQt+CDQg3/
tl3Ujuj2T/b2g6eszo0f6haHpG0Mxuu2MHjk2MhIK9+WkC0BCp7l03V5Roa4wCH/I49trobGczSE
Hu4TWDUkSCJeNar0Ry+XjmBKMYoAIIbDwxG5Mtu4idtI+6vCOfryq6r0b1VDa8Ry8ivjDULF+ZNg
gdTo236wR7hU8o3XAnybi1pmU0hQkldtAdaSzVGkGXrT3U+ftQdTvF3KJ0CN0TH4OIYc5zSxR7Zv
nFaVp0JekDnw5CRtbbSHzJY2vBL4sWTNhqeoTEje1Tozjvvc7selwhIcpDpg+QCWVmDnmdyUrZ0P
D7o0RMpHPHf6TiKT1O6r74VzUhjYsWYiB7KMGovdtllgSrzmnpq+d8151xSYCElD0AwfwJ/gKCvU
ZqTfrEvxjghMIRk5ylguJkV+Bs6VUu9aznZ4zWqzHqnVk22z7t7g/b7CAAOyCOhXCTT9LsWhbn01
GtuukNLwtvh9ZB0wiZqb4b4OcuIN/wFLGB/zwcnI1rhdMoVoCfOebDNQp4buaoqz2o0UinvvRhgg
Ba3Xrg2iFGMySizjpQQqBGDAF+Gg+cJfwhF0hKTi8jIyV6GQ4l/2hOtxv5tgmeR8IV9XCia/w0o7
FmT5a0Tq5LM1gAUsBjP1aD/kcOJzJQ4mu16Ftm8bqTssBA5K/gVVgwV6/UsTEvx25QkeBOax8E94
mv/+CQ1J7VgBJB+qxcGwj+KiHJyiwA8CFnIa5SLcO0gnt47t2iDUE1vEo5JfoLwrgeyl7ZyRM9Ww
QzshSywtFV8864t3CaFGoCMOD4c/PLQirwsdab6bYe+Jsh2Sq63JNZPPZoF+QoVUhOaUGMHqj6Tr
NcRlMTqpfsK5+Ri+JfsQtIBpNhbEvJMTo/pvOjw5rITGIpAu29QrN6k8wcQ8IlfjEkgPQGQ36Wz7
Buo0YTVjuzCEgtOtymnyzqnES0omKwx02xP/4G10wAcqydiZfJpoQakxOH2lJf74Z4w/F0qR4qzx
DpyGqamZSuxCNS+Z4Y2gbv/n7q0L/pxOzRTSYPU6dhb4+H8ZVSGY+lYwjubutGjjxoH988CJ2YPY
REoUqATenIz1FhcuHAoxk+gpdDTBV3orIJjVuHMLl6vlSuJGVS4vuKwB5wu/aFuKTAhROTdOVqM5
B2XwypN2d/Vsk9ZKBiCtUIpRcG4RMMFE70YQPtEj63Mk0PRm1OpFM2kOaJnDJ/1vEBsd7ENgjIwh
x1bx8tWJDZjSfUkXHc7wdTnKZazvOnclsZwSKMEh2Wyon1416rAZiype33ZS6LWjWpSTy0bdXwG2
3VMati2ZRArQJSdigKFpnllZwwaYdPFYzWip53yYdTZ4xpWiWeBoufU9n7SfGWnPOI4v+H4OlSQI
YajHP+q3MBysQTTqQUzWn435F0BKL2o1K8s+dKjYuccgyyMImf7bOWHqx0lEl8j4Vhld/iF8rmZ4
1mXYKRnfM5D48f4Ux0P8MRLOdfEdYmNsj4xdgHDBTieyj4xZPIEphTvzXILrb6W1v0ons4Ji0DTJ
T7BRW4lGJSrhsXZzMbzQQp81HTs9OCKJRX2tJkfODXxuRZTAOTwYYjNAKLH1aIjMrMsQnfnoxoPP
d+crkpjhsScsWwfbB/AoqX4PyOU8PumpDRg4OjAnC9SDnSqFewwdROEXKbVqqPw8P/ppLMH/inbK
M5PDlWYUGi6O2qzgEuHNtrXbsHysUYmArwqjQdLMqJMzR4sY2WzIQOtB3LO9T8BL4D329arfJBrb
Yv1TZJ1oYRlM8fcOCp1pMAfNxyR20OXWYLZjOs4k9edv3QgdzfjAOqROq0vs4/JzPqjzBdLSJbQS
RpMsjokfoE67lMLE6PrN59k4XMLfGI3tSsFMZ/jrhLqL81EXDqeGD+54fEEh0l1F3nc43z4cYwt2
rCwZZiFC1uHm3JMA7heY0KLDm+VJ9NhHzFt2eX+3CwAgIUxAN3mOkWama1+cSaVR8gTuBDz348Jt
QMIZJezAbBo53/3lsNsg7MfDPz43gDbcjOeVBH+9wvcdlS6Q+bl6ldN1L+xsCzG1kIL4NRPeULez
ZdtcGyGs/SKIxy2fG0W1bekj5PNXacb9uaATDhPnMG1oE3AmQ19F4tw2TvK2Dbq/klhZIHC2ijMA
UQf0c/1203umxPR+Spzu7ucoupD8BMurwYgNJMzOPge0ji7NWlmzh0dqmTeEMo3jI/estRzP+U77
dn11pv30jX2e1OS251ciJKed+WIPU1Gcsx/0mIYmnq857k64WLQ/b3EugNwvDkkJX4/ELdv7PJFx
tGSU7GTrBvX02pruIIqyd7bLkb+1d7GXJVFB1jHDieOPRqBtGQFHd9zReKt6AlD8/hK2TMJazvtD
DUvlEItp7ijZMxPCqmrPPtw2tOJxOcjz+IdTZWngB3ikHIEib+KciEpatjNn7Lm0vwCPN4M+wpff
ATlhCVhztwuCu/5EFUb5G1ItlwnIJFPVi6yKEm+4m6UqCsAudobYX+ynFtLf1B70LqCurmnYiR31
x+piT2WhqV3enlHOaqcexEh5x7SRewg5wEBcZzGfaL+nBAxMlXp+Vc/Ljn/bd/pzQdATBVPawNk8
xMmrhmeiO00msqgxebXhPVihAWX2Iskrb6d76OEtozBA5TiOmjh6MZhjfsAQSihFfaBkIPO5noyh
gk8xBdGaSjy2EWoJsX0SSmxSpAbGyn0ZhV72OhaUmecvNmMi6mzr3GL2+K0BJQr2ijvfNAAiVQot
PzvFeik+7ALd+0ngYfxaUjgv4+vOHDH8/GxCEVDunPR8TTEmH3SBrY1WI7HUsQ0otSARxCtDEXNR
/j5WDDOPUnLqpQx9Fhu5fYqeuOzCcOwuILufa0iA1+Ag44IvGU24qUUMSGJzulDiYLm4KhOv9+66
Owa+yklEOKvjk+ivrsT8ffVh4t6CaytjJmjVg8rWs6Gv1aMZhV7D+3cW9VLNnBE0+Q6dAaPdu8ve
DlBkGe0VOkqUdda8mAZHWx0mraGO83W78ORR1RZhvKwXyqkjIyFYsJh5nWiv+/q8Nkp0uYA4uu5e
m90hXhI0qro+VPPoRWU/nJgkT9VIpYo1gXduBd7Ru5/djR+chF7b41iloNOStkT41u1pybSw+5S3
vBfJL3jpCnjxSnFc20Wf437j7YPO5UJCCOwgcoO+33GTIMbjeXjhESIlSi/+0Nq0/Tplit0t40L2
dsTPDnVv3tkcM8UQmOZIlVv1rPrPJ/KukDvdwDwRpnrMy1lQ04GJAqSs/5cEZ8rWRM6lOjJFXhFu
PMWFU9MZVRet8YUVvEslz6ajpRaIC//Au1jj7BQ3fJgap3jYrSzWl3rpBcT0jfpVD0UHXpn2p5wE
GPAIoKdr24DBtZ7YMAi6NeD+ABLwQuwYHzvHS/TWcxCQaFuda8GVN66NUrXXCSEhQXFjc/PqZXsN
rEtCUDcHla7CqvsM9aLRp6lR0ZCkRejtv8EMPZD7+DTBpt5UJu76tIwZqw1egeJl1a5lzJatQXRu
gWbwbYHCmapnVO9Ia0d3PgJyfia+RxrFQbuIjmuaGbtNR1dFTg3yFxlx2d+AytnCRALVsBd4ATU3
Fy/W3wltXyCAG4yfdXhgRXQCYICSxd6tYhpjXmxhHYTjGgpuO6CGRgnVhuYz3/wR4hMJ6LLa6cD+
FTspBDGVRWcPUCGNeY7lsM2lyMXZ+wqQ5yQsdZenySjxnesG1JQqNWatHCbn+OtQ/JAfBNXgR2FA
6zNS4rtaPGZDqxY2jp4BL4hY0M9pgmZPXgxasUa1ZcW8ZXErP1RF/KJ3NZsuJePoG2jOr4yVVvo0
YrwW3OZ0Ie10DSV9IbMuDbjEoLUqiPysBDeDoZckbIA/vhCulq8QXgmOxT9jxOizehV5hngGCNgb
MkgEQmr2RX5J4AncjP6SLLLAXxCF8c7zyu+OZtCq9gfHg4vDriNTFsys3oD1lgT0SnnraVA01RCs
70XcYamSC/8YCWd8L5xLUIdIW7nOYRD8eUhbXuDWwvN06HQqJdp6g8kmSEG0x4Gy7W9pt70u1RfJ
lOc3CYhLjHvbnsN/kyKhcnPa73bkIbcIzaPHnpe7A8KhgyCyjRu6jAnRqX9njiLfdbTOV0D1v+7a
5d1JOv96PH9m1ZOMP+FIwGi1LjeUwrd9wni73y+7WjqoeSpogZCNEW6/ItmW/jK+NCGz8+xDvSaT
l8rLmPdhoJsWqerGYgcGO7cQ5CapUrvZa3d+m03BAxOPAIZMd4LA7QcBZQrtOGhJ3dAMPwN1AjyV
7k+7RUHm2Rs8pXIejHyEonHeOjwo3Yn0FvqMZyERu4IyB2Yc95C1/R95WTYPKWNJZWXhj7LkzO8b
p6dGYXfzpanJGyO2O92Il9xa28DAxq8ahfdS1SXaz+gQFrDnk1h68y6GUF2fK65gSKqD4ADDh5tq
xPw9xBSXl/nEKjdFzAJ7w1mth5XI44pgf9cCB0zUl0oYzQPs0RUauixLNwuGkpkFq3ox90KefHj9
R+gQ437RDCTFAspf4tOCEN7qLNmusOA6RahKTLZXYuXlqjJGpI1HUs9w9dHAxPSyzVqejYT5/L1N
rHZBtcdThq4uvuCA0X9Y5Tne7MP+jgUwvSpQLFYcrxrtFANnUxDyRkPgOx+vKE/xFIuxnMWs5yRU
3cLgVQ3lL+SsTw7/sHkqeJnNum1QJdE3EUlGqEC7vISNc+uD8gPmA6smF35AyBXTpZbGiVhrNA2+
eorlPGkQp46n2pWuTo2dwCKJ5cGJXFFzkIaEQgFhOCX/g3uhzn9PQ5UzMm9UQE4XVHN3r2hm0Uq5
ryV/D0REodJomCjIdfXwq2o5T4PW04PO4iu9f0qMY62zcTCu+1NpEt8oUL5XTna/QTDd4gPdX4PE
OfkiptsFLqi97hk66AG5pMpzCn8Fq/9uUah8ebJqn/guIc053oXtW+O+WvZvMwxYi9afXyAdxicf
MK5rmKOAU7Ze40STBhKNFfyjNESxDPPuLMknh5SipPHTaU+VkR/NdHV+HxchJ4c6kSZkKIXaRdSb
1zDy6DpfgXYX0LkAAiR6B51gxn3a21gFdAaWnkMqz2J4/P2it6YKQep+YNfH3skKvYkwZ8JZDOCC
oeHQ30kLhvHq2lVCfSO1eF0otCpWhv/CNQDTRBZbMJARIvsD6sFgUt9gMRflEan2Nwx1BTE68CBN
RMg3pwkT1QHOcY+BUdqoczSNDc5PafE3yt/9w6xtT/PeqOnoxRkCLaUR7fmwBEZbIxlGtrwJPFMv
D7RfVTpRCps/JBcXR96o03hyAMp6hzfAxYIeiY1/A+VpZ9KBKhq82YHVkgaFH4dclZW3UA8T3YIq
X7r4JJk0lC8XC4QUoPfUeh77Z53xObvig8y8JetSSrzlQReOAZON9rKHhw10g8/agHN1b4axpOCM
iyChKcU2hCq6SZ2P02MicnydvYzV7FsjbSc7bw6pFTdVSXp3LJxSeXBjuMHngQgTsUWEqaLuMU3Q
uphF6XTgvaykjqDilGkoR31Z52sMhOlcOka0l2ikDGZbvESve15IXLl5Ad+kDqmm4TVF6fVoNk4N
WcO4VFAEaVdSKJfJiij4a8g4djurSyVDo3JZx8gfOCM4oc9IC021P7OMePGcUUNolpR2Y8nH9hpe
bI5VYFXlrrmLEHW6xbaaW2lZBpTndXNgnkJk1H7ny9ucfCZ6TPr0F9jxg9gGeF0ycwknenQ4i5TF
A20a5miqOWG3bnYu7IlhWNVBGU22CtVJQ4X2sdnk7UG+v6FDxyAUpsxFgIbgfd9zsW4boNcLC2NH
VjUC4iSAchgfW9AH86kDgOhLl1o/+ecqVI4l/opUkYCnk4LK570yeRM0Xfcxh17lwa11cksIfoqt
1kvHgprkSaomGKO22pNZyrVY5xngfj6cR/ApCt+DEdQlMaAVe6Zn2GiAF2wuXw+oJPHHjolHokVP
EuEdkiwz32h04NDkQIOpiCLIBzGbHfvDnh2F2fpH9LOBaAjifMKJLIpU4qXfYwBak/1EjiOfYyl+
/nokoOAgaFcxhctH+hkPybljlLtauC3WLpf7gvFzGPC9h4So5AwIryrDT7g3fGJD8KQty6Khmjve
udvLmZFDWqApukGMdwuXZksXzigccuIqHKVkLJ78n5kk+lvO37dyMIiskNAzzYlaZNsHqsk6mNgZ
5gN9HSCB8GAgg0a6+LmI2j0Fg3wvQpnVSjHS6r+5PfS6pLJpHm3mEEYtbH+57EwGgccBODSDzKhE
oLnEVWnKpaFWqyDP0yMD5/k5dyTdujHPGPhcZgQSEltTuQMJK5kg0q5MLdIlGbaeKDP0Pb8u8DOw
/N+mncT2249HFYB7Hgp5sEgPvDotIXekbnjCDlpizhnNlBBzl9MDJP4XkS48JYHF7mSqfbcTuygC
zW9R9nZPBgyTeRGxpvHaYL0kDQvjk2RMoivgK5jBC8niiD8WtaCRQQXutdJq6NRti5M4vr348Q4m
rCbiScoELfBHhebgh6qmsMk2fjzilpNtdbFwCCPdisIbNPnwKjCTf5CCIvnrjD8VLFbGbK+MrjR4
r6OV8nR3SRmeVhLUcPEfdIToMxnHa9kF7i2WLEAJBRcfuuYEYMPUYK2XBepb9A79DERZDeZhV6L3
ybjt3/kD+1EM586Hp3+GFqM058YliN/+vzX8vbB+IfgtPVneQ/XROP+k1HgJYf1dISOJv2zdF8AQ
UG48NkSkeDP+Wgf0n0SjINV7fueSktGiMacF2Q04X1Csd4jGXxbO678PKd71SyyX3GdLVqq2o1Wy
7fsE6gHF2g5SzbJsaf0iU8ddiAGmWxHMjQan0pQe33Y+n19JVTrOoFI6Q9kbIWADrx+YmKXxXg6k
ZzenaKEkIQ6mp8w3B220nhhslFF0sUZPyyz3aS/xgPdRPuzdnUDpRtPI5MOe8kwGvCt4Sj+jn2vU
TF2xA1gRCJqrsB/ikDFuKlgTaO3cTCvKRalOreuF6qsL6PlZaNxifycyj+BkbC6QZC+a9IIgQY+4
XO3njudi73VTbxBHR+PCbeIdsi1hNnSbhPZrKIS3qH2JdnYyIAmpnFuKAHlxUOlsXoFzRqKts2Px
AFYwRV4zfUnfU69CLgK2OzBhWUbJUYEV5H8/BuBpV8e7HpuIUPqlswYG2wR01FX5zOp35Tw3tCIt
LcHQslx/Hr2VwATq1i6XYqo4u0g8MwkwbCD4OuwuD+NgfKQW6+APTWQiZmo0ZbH61+rbs6SPh9lz
ZRZSNvD04oSO5TQxfqUT7SuQERJ1exLpmyQiwEz6CfIaBl0tNWnWD9QsE42W/x0DLid0dc8G0G1Y
h4gJr38YxxpSpySuub+c52dqVMKJMlChUTDcEDrdMdTKtCf4QvOR+JfOUm4f7naA5BXb9DO//EeX
UN86Ivs9OHck8s8BU+ag8E0uhQ8lodWp4tmA7Nb8ll7WbSByl1NKOci52/QWDAG9kpEtE8S/xRXy
T6K65zCM4Ebw+AUFq2piqEcBV1HN4+kHbOASXL5rZeiZ+1Ei4DrHlt1lPENOM14F83TnnIu6U18r
r8amgm1lgqQ8vpfEPwsGC2nr9r7LA2qVLDS81WjAbM3Fluh1wgMKZA43eeRy1CpiE+Y6cJt3lDvI
s3kqCYF/iEdoZ/FLMs/7zZWTWJ8ir0j0Y0Ory3qoG9LDzc4Q5/woPjamOHcNx1NLjNBih27UVFPo
dKuDZXMw6LhtMNbB5Td/fcVW3BBnZqX2hT6AoysE1rf5oT/eFrUwzcV/aOwGtpsgezlm2FAuXIxB
JVYzXGD6e9wxZQUGdD2IVn5gXuVepTNoKRUOziS8JHAkCZs3/MShR/M+DA0JA+RZejD/+AVHsFCv
i5Q2yS+ghiwQMW6fknu9eQD0Eu8MLYXZP8hMRxHw8yLURy9EqAThj2SUV9fLABlHKUKGN++qHQCA
FL0QB3Fkzqycm18ZbQThDvIhxvwrrLQpCt+hbEUVfZZROtsih13kNiFB8r5/0A61XSLjdbyt9x31
EmRE7C00+hqJsWOil/ckBn5LT0OBiIiRC2wG1YBR/si7lgJkS57pvhiwKAMZBJvVHlwoHDkwhgvx
Vf99Lt5Bw3m5hv6UuxPyU5G9VB2QjrQ+1yXLX4CGSQJfLg8y0dHiBme0F8y89HZDJgGXmzpQm3yI
ihJ0dZk74SqkniFjw4PJcTe1PJLTiNVR4vajqNOvGjrZIB9iuCJJzJjSr+rOS7CCDwa4gOl5LzP1
b1P3Ckc7Q+Gkjy07mr6PE1tqUl2/sEXqDAcITlqfVb4jYu7k/r+sEtIVidFHd8AV2yKjIZat5bh5
43wK3M8sWR11GltBdd9CCjT1rd3L/+qbuMzcJgqpe8XqDNNvsWguKhhegsIEy9tA+XkyhQrmAomk
o51xr8YUHUMBn8X4URiA8qj+jD3mjCDn2iaYPl8xuUMxmNnNhjJJ+P95V0GdUh5NTlDA1iO43hBM
vc1qnZONefzUlvtYB0U3wMp2LZpuHJhjbAEOXgJuNctDsIIYqGl7w0CFYrZ/KTtvdFboeGEbMabl
kmSHRojikgZLiUeUo9Xj3M9Rt2K9O6P6OGBdAz6G7SgKHXajSHeBirW9MB/aJKuh+GDphme5kP24
W6DA+YIv356Evlf2ZhjpcmZitkCjFkAtLvhVms1j2HkFYfjhy985/QzqcKHzdHI2S7PNQTLwjreF
x4v1xG98/TqV2KgoQ3RAHfKVDD5wg9ieRLP2VQgyNzQPQL5e6a5sqUcGps2u7F8xburFWHcR3X2n
G9V8hWLvqpBBHiyXdjroX9Kes0u/RIbA8i/t/2iPkYDIDsnD58LUtDn8scTKsindu+aJu07cXwK8
yyuAWGs7xr/ih61A90lLXZsvPJ1KeMyNEQ/yDo96/tukrvNChURr7Cqgh0Bqiwx9JIzNlubte1Ol
pBH4flnGzV8jKTj/H2foAIbpYmyWBHh7ZLMExUHce8EgSXKa9Zmwdc3AY5cID3APsaNswW1PGuy1
tvBxiIuEdAr5PPDSuGEV4hOaIWOhA+YFLiE7PMw7bCOxVSNc7WqjTpv3AYp7XM0k4l3OMOLkT9Bo
XShlXZuA8Mvr6zav0jOYaS4CNBtO+yAG4mMkCC8kBU1TNcrVSWFqmYKv9qnvzDlKb+CMKaPsaUHs
xH3DshhUsYHvIMYN+mbmfU3T2g2F+rSz6Krif2wNLwkSFm0QqHj2xL1U2CXcPRUBtK+eOco6Ixxi
dNmazGQSIFFPArRB1Yes1W8IsclHo4AvVsFjLYsdQTEE6qqXsmobjaf5AWgznJ54xVJUBTmBgeAw
b/AdOEJfI9exxgy8d4ZTw+P3xPoGuhFULRJaHe/Au6xGCa07c7hLBz7GNwiYNSfDwreE3gquvqY9
vSyoyOyGJ9yU4Wz/xwfGsMjBM2RBrNnCBBmeh+gN9+rOqKtAcP1QPvPXk89tY33vORWEYwQk3pJa
2g6Fs2hZ5qN9TE5NxQA3pVfiqCa6Gcf8iKtEG2AXudn3ZFAfK8GCmRpi+q8nnDHjp3lsE9aLaJin
Btt1iY9wBtyo3Z1CpFQ44hWqZTvJ5hSqFQuwkquzpVgFe3qodwY7wPSzPQtmHv9ZbnwEEMkdCNl+
pGGvwUcwK1pMTnKtGG8oz1UrWZVYw0WiF7oAiBzhaMTIHTCxxwOnRnnNqDEMTT5k6fteEa8h/aZn
HmSpeFcks2DM2+8JUn/zlnAsDss0ijmAb2q8Zo/jF+KoUO7TDI/IDTPIs8hcM+gxgwUEQ3q7aCkF
nxpG3wpkPceaCALnOBJV9xXc2FuSwZOvU62JEdv3OHoOxpBRH6hlpr+mnw2H+9ukV5ggOP4DcDSp
Z+8xCDvK9At/wIubktdEM/3MLR5nI6VSAV8G1zkkcXfQJtjdE9bwRfZMJIV8Vu2L/Pvt1ShNrUCn
ckoIq1eVkaU/l2G88oAaPEpky+TcWToMXb4WoN0GWoisoA//H2t+j10LNsj7iUZJQlc6HbFd1MqD
xuD2j0Q58WnszZCA25sTMZ1jCDiZ9EWX0tlqUHSKV2ammCrRdJ9I+kbqoI0T/FlXHzFYflvwATvA
FmHoq5+2TmMf
`pragma protect end_protected
