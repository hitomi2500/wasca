// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aWVrFeydVbRA78P/XktACLkKkHw6w2PG0dkibtpH1+PZNWruXI1EpKFaocFm2MLuyniKlj0MR/3f
fOkJKWWGjRWV5EVtF5VtjXUFA1WTHIE40lyqUhZ76gKnMfhrXUcmeb5kNCMQtE3CWyok5ovOgeBc
SVrl3vlf9T6RHqpcjRSii63yc8zhU50kD+Ste+VGEPQv5kMxnBOTlOPmOLNBiLXQojbfQ7BgQwGP
srzyHUoDlrFng7UkuGHdJORkHCg8ECnIvTm3ya706V89XR5pwONQeEXZ2vNxNoj3u7NTG+GphoyL
2gVxkdG6GFtk+S6Lhw4Yp6fs5F9k7epdDTZMog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sFMBy2QMViIO/S4wMcF0lsEmucj4FbfHdG0cXyF3lDyEVaar9DQjtl/jpMfJiZ/uHn8VgwiUEjD/
5vTPs3yTBuwA7VIxjJ7/J259V4OOEdXFmTN7cR197ApUllCjWX9iUqf5Im9TdGibinTjeSlYtzX8
IZLm02/wrKxSTNFlignbTv/bDnkiiBD94Tgm1DY8ORdbxJR/dSXwhop9e/UmnhzXgUyrs5cCxkQn
6a7pFCLYESD6splU3eiu2te80HOYDu6TS3mck0rG1ewUqq3afNxa32whKX/giB5ndwN8y81OrGsj
8VwMdSzJlE1wglaJnJ5iOGIw9o9zKP9/bocXU6pkPPMSnO8alYwpmaF54DQDzlWjChiIwFxBSM3s
hHk6D+70RkwIQ9Su8GguuLzOW3Db9fk1nd646v7s3/5JgPP14ugnj2Hb2XvnMZE/+EOxZ/23b/9R
CKwkwRkoJh/SNyBnqVb7j4/wWfQcr20eXYEKMgHnzkCtk2yG/3IFIVTZFjjTEfoIalVQhNzMmtTw
B+YjPyRnHvQX2jngHx/7IrUUfkH+bmA2LQ9fEWqetJocuqIg3w3PmGLBKAsMzlagdBNYyGOw7eE6
rdLP/vg59E1Lk2M/Znd8Wv1+1patp+i4wywBiYdR1l42IPac60HlBuDmnBK+5gqGnVVxlHZINrUI
Kcm4f7zKfxeX9l4GlQY4IikQGJHDzJTanjESf787roAbyRPG/OGOGq6IxewkM5VeppwHf9rxpZuh
8OlDNz4BazYEvyH8ifGq8R61Yuj+KWh67SIQmHBHJElQvPgS5ypbwqptawuKckpw7Kz4jW6RhDOl
6WjhDy02lp+IFJY4WV4ducoLQpjUl7k/x4KSoK/WE3hbAb3rB+6G3Pp3+tk6S1y/Mo9tbtDbX2Is
iKmrq2ezZvazY8ZtgZ38+8v7T57QrLJe2Hl/OX4tevpQYwAbAki1B8oEYa1T+wzCzmi9hLFOrVht
RihZok283+aLunt2HKN0EDvjb5cxhzfd0KGp2B4PAF9kWL9fJBwbJNcnc7A+IbzB7zHTCJtGbzV2
CGDXJjiTa8X5hI93UUCZUB41HexAlnFimACerfofuUyAvMkRzJkZNg9d1VIf35ipq+mUMkZJOxfw
bfSHcwQu5uoqnDqg6r7EDFYZn9+9dCQYejqi58AvBFnWwgA1kf9QyJsa0P0OQirfjjqjV/MEm4fv
UYK27w140Zy03hX4L8yYSU61TJrTIE8tLjU8IoisI6QK/CGB4hxLlqSy+tSajqUZ5Csb2Cxjw6gx
FrVZ1sJzq8rLhXwVnmdYJtbEyqt9sotr4WyeZpSvzxMEvxjfd5ChEqnE9tb66hV7Fi9wticvPL0a
Q/Zb8YgfYfussuzWrMCyw5mPBE3vLh8Q5o16u9bBL8IKbljvoVvMpipBeLXzLtc3Cq9hkWH2D7Bc
owKmm3sdhgfEqgRgXh2XVgpegABRHtSlxsbOwCXQJbDSrHfrT7/pzibG4bY3R1Eec+CH6kse4eDc
ewn5etuGxbfxZH2le475pE3szZSEdq75Zx9nRNg673zJsePP3JrD8e6p4u6Zil1Rsd6Sn9WUbcEB
WDP7F2fhP/1WhqYUAElg/m+jjIKYfp9JjpHIxStpTQ8n94rY+VOCioobNfqTu/m9ax9ZVH2cXp7O
9V4ShAigw+MpVa4guUu9qGLtolRXGf3I9zBu6uL+eELir5Hp9ztgiFCSka2fV8vKqdO0crcQF/ZQ
vdmmaOsKjV0vGh9g804mvu4q0WjIrhasaxlcwajQUz9OEU/xgAt0elBYnfl1ABxH6Vi8ToVI+one
aBEMhFYLoBE5k9vb/uunZjXYSdDxUnFmNyOaUF4gIDouEfQACv1pgQND1PSdzOCrzx+h4D2v8W0P
ZtakVnETSaiTa6Q2q85sZFBpwZ1UA6lwshxH5jeXv5zZGL3WOTAc5hjlNFcH4xm3iwyMezi5ygdD
GAF+OiACR71tlKVe6VKSDGqYbb0ZQzWZ274GuhhgUDF+ADV2rxgYnq2B7fpGpt47YqYJ5YjyieDt
njBpu6mDYcLZrC89oKfd01tNTN6c4NtSGq1pxukcPHHDob4GOcY3l56BUvtAoy6GjZY/UcJDf12M
ZJgdXNMhDYZ8Y+ufRbqJqL2riyP6c3CBNIE6EeDYoFooL3mLP8+frT25aDdSzYuAVqpC4omauKTV
njCa1108pbXDDZLf4kVvnRe+g9O0SkM8C553p+tibIiasz+7P5mJs034E1+uaiHbBslFtfZcA1rh
lMxx3aU/QXJh1hw+HWn7T8ARhC6fu/vipbDs/6KEIPi4yJoLJbL3hncjFrxEqkCo5pRMgsdmIY3h
M3DcqzY76NW1MFUD+Zga8i20wvA5Z7+cRscokMxt/iK+tELg5lfSKP9VTTudKDe3JBY17a7JD8IV
8m9j5uooxdfPnsOQJKdyCdkM/SQdHJKaNYMMIARDTVw8fnsuH2Cu7N6nDq1+/tLqDJwVeO4IFn6d
YXHkx7thQCq20y62lI8qoEJ25FIa79pji8yWMUxkcRZxyzk84Pfn+1CNO0+s1AJ7pQR7xCovwEXL
GWabnhFDIq9NhIhkkrxa8MrlNeSziBxo8mzDkOVhGYxkFVdSuKtpIm7uR6XgL/9YonkHNYl6SI/w
BEkYbFcoElNvM1ZYN4ZDVvSfIe7fHPvq8jSwCkoXb8iMd5LQTfBUFyaZcRzegPAwRhBHS1c3zChw
S82IwsFwJSODJayHRL+5mN1Rp9lyimFKOLOoqz8SJ9ZVcQtC1YhgWGEIVviPVuFI96fjgkf9QAow
jGwj9eKIu9ghgg5kLeU/mSXRKpGo+RhB9u98M1GctqjK4LC1NydIhBfx/4nDoIFeVfJfF1LcRdmh
VW2//IfHIvyuEay7Q0mydYJxmMJz1syd79RF42iQUhww6VIL1QDBa0SpqOS/YlSPAAgB56x7zYPe
FWK5+h4DpV9B0f5dlrqONoRHg5K03ifsGxMHgrc+rD+uMO1N/gFc+7F+lOBUJQ6bUhJV/GHmXPgB
UiczDd5GAZM2SH8fecAO9CRL49+z/05PQGVMAjOm9AydAnevJTmMDXO6t8v5scbwJmbIR3YOHeIU
pKgdUoFD7J/a7pUs//sEow0LPqHE8MmQ5l2DPqXUtFTyO0ZAkt+dJWyT9CufZh0PBSCZmff5jmtz
AjUp+wVpeMm1ewN8jeYwBO3PC3hMraGyZ1HTn1Xeyfb/z8EXjMhI+M19FnHHu1GhmMGBEdXC8puL
1wCprw1wfsfcYhQrWQrawIVg4H3a/5dvWUy49IbGLGahSoVSv53fK8pl7pl9nRVoYxiF3YONXIFu
i+Yzz8ANxPXeQY94bQxR3AJ0zp5Vr5OQTPj2gvEWQ0Zz+ceV9rwbjLMVKrla7G9oL7a9vjhxZrqE
V/IfIv31gChdMjM/e26dvHBZiRb/H5zaA8VgpK4i2tSpIBZ4Xisn4GIxRl1YAwEmQcYoKy9/edAg
Mlhi5BoppdMFPUpTCw35oLnNsxo27LoQzdcZeTMMoEes4Cu1tHJdNnhAebkuBocK+DJjGic7+6ET
Ae1Ymm69VE1Iiz+7nrfe70BNrJBKlXmgCrCsZ5iqEXnY41qEmIcWuQ+fES/jPg/J0nJqHE3Pw5aE
Rmco4z7u8pignEy+9+P+rxo2a8bJYaUlaphsxhy+1TVmqjCKXlSQxTOCT61hc89/jLa8ks2tK1PQ
7WboD/eK5h8QseQ+HCNrrMpfnzXYcuYAZ1sznH6guTyUBR6l4yDXnqez+1wtVKIesH7K+0KOcDG2
6VjJLxMqJqt2Pc3IFWP+gZsR9WxmlZGx/f1KHrZP6Ox6EHF9bdeD1STyK4FQWZgeh5gXC6y7Ylh/
PrLld7OrUAqX2yGFru69NXcokSpKtX0BhYFysH06nVY74BexRRId/V0R9JjuH4cvnD+hoNleel7G
FAtpiHVHZfIMNl9eQpEW1DmG7mPj2Sh5+ckPDOR65nykaSJ8bvsFh1R5WYZ+lTGTBEQeJ7XU5M9r
yDwb+UDelqw/0fp3A+RURiaoV/GsrPf7RQUUuc/dAu5OfW/JjN/pDBdw34GXDg0FIEVffS3Ymwl9
Q7bFFGP+7qEe2kxybrV0GK1sp7G2IEJmFTYzpXB+MmLA5sL+ipKSaflZ/zTwIYblDY15h9jowz0D
JIVG6A6Z3ObANyWzhkGi5fH58SDBKXRG+tS0zdUaNgHX5FEuKm5Yz0pmJ4CCgmKwH4t4Uu7j9nKe
djws6z6DwojitwePE1qkx6TppoD8+cVUGUsu3t02ALy1h2q0s0vFQYfGbriZ+qR1R21wOBH30uIm
KxCgVG2kfyFsBbU/bhQuTO/aseJHFshaB67Uk4PvhfjxVwMTaWmfM7c6kgJVrhc+XgCT9uUyBYf1
LoHaZfQYZVcmxvFAHQZeTPRRGtr4rvUfC4al951PvxfSEF3xNKJPTHeVTCIaXPjQtaIU80KiPOO2
O7S15wZIDyTh3NLN6z52bGdSI1CAW4ZnB/gtzqMHrr+weWmZ2Xb4J9uQALLx1cyE7xJedK0K/td/
hee11+3cg1XGQOsNQ3D5ma2nHRfTngRBbzDaGvlphvvWXpeO2+5I8xdM7mDKdegxAS4gPSKdFHVN
I+xPkKN2yFluAeEi/wcujYOprVW47JPY5Oca6HtI5rQq6XWzcKeX/7ByCho5AG4IzmX4L84l9KQD
DQwDFHjT/nnMGg0kSXK5P09FzASHYa9KVhkYNPpwz88GhiSF7nUEOmma7OnMQ6LzEMNh+I1KkHGd
XO9MCtjY5RY4HrOJpx2MUumvJW9cCvz9FV+9D/KlTQqEY/Iq6jkMM23+RdcNud+CntdKSTeTabZa
GtcInrpLKxkT+5EV+EOhQB/Cs+rai1uCswZU5gWcNylXpjNlRm7pKoOuqytfl89wteEI7e0q3E2W
0beCkKAgd+4P3yWM9RkgScJooOQMjykr0pi90oYx+dO1cxK22ddFEjLlBOdGzlLe7INVAz7txkrM
pL+3QfsTuCOOhpq+UOcNcFm/+7DmWGF+jq68Wt9pmbH9qlvqiaNhbR6iSh5dwjGWOJLSPurKYZWu
R2/a7j4MgIfCpZNDs2gyq3V0DDlNDOjBacR+07WIp0UnfA1qES7SYivD1yRuLcYbBUpQlrPDa5x9
x95qghesaPVVz3XPqxnU9y+5QZkI6UljvC4P+YQt8+fsZCbPDR8RczMvpu+SN0nJKtcHFK2UVbfR
hgtQgAR0s6L8TJXtkFjCtSr5U6GH3TaYFjivykzfXSMT8L/srqmvq42A8XlMLuKVgtFPGuVJkb+R
9UebR1Ts83qDWDXOk3D8vLLLx+8p+ZdHB5HEZ5AmIxxYGqAJJqO470PdZBkZLg+mnUIL5fXRhtmg
aCVfLjpAXMZ9UK7KvvzrCoP8rjZHTdUAoTDEjee2Z5RyyyGRu8PE6DLsdfhsd5mv5AaxcncwZJ6f
UTbqDziqA/r+Pf5KR31519hhZj2XsgbIo21e2R3sf6BWwooKM4LQj2j35W8BQmcBnEk5HelclJUr
xoiHeKVktPZuqsfJPe9bICh+rzHR+koZLkLS4YZvNN3OjDe6VBWPcYEYmE+X+OGLJVskvgm6Xaro
JpjFo0SOICvz0s2rpvc8H7RdI7LtHj0LU2XW0EljqICtUq6EwOqMte/0agiauEN4jOZWvMPKI/cz
tg+MIRbvujG0NN+OKiS6UgUp6u7KXsTbGwYjxnlscDcV4E9SGzZB8lkWF6lADU1fYFrseyOBHJjP
qI9IFH9HLLmMCdXgkrfqKOXOkfQAelUEeg0V6771SvIJDAXHOkR8JkS3LS8Ge2ExMnUEOet4yFt9
3/pnko/xbthBwbD0fXhTOHa6iUfmhXeSahwDxmtjgc+KMpyK10hFMkpdFnMukvUkniOkzqIM9aL5
sNhFcsOSgnpBWAMellFEu16xcupbXyTIl5EHdbiKc4JO0icZaGR4o9Hmad99S6M6jF5MvzSR3nvc
nb6xixyAwPYIX1getP1XBit5nL2zPuQ7V1eeAwKmeXfeFYNQJkx6UZV1CTLa2pzVN0O4JUDPcdhq
4KLd/+FPXIXxseEWdTtl6Pz3ZkxNKNXuS3JgXUsHZrVDabqFUXARcIc6YKxpk1M+OSj4NISXaPl6
xmaX0a9gIUmQx6VyllbMiKocYaltWK93kJ7l8en20U9KSxhup+3X9/S7CL3REjwrsp6DDQ8G2BGs
fHI+AbHvC8b6GZT6VWiH9wN1sI5tydUp+Bm8buShkNU3Ikebj6FHKe5DN9fk61v06CWf1KwHZllm
0dU1+udLPwzouymXcs9kxMhhTT922Ko0WtpPCPj+zpaUG8VNQiDMbA6eQ3rveTKhsCPVT36lXPj/
DqCqro0ropT1G/g7DAgzy7dl+OEOQCiTaxdrcMm0Yf8eYTN/4qKGGMaEUOuInPNlTd3O6JQwngaD
OUhhkIXqsM+JasskcS6OVj1OzfLUtFcAS0KXyzIAv6IDUUDGwMwraQnmvZ6YHpEg57p/0YYIYhz8
4sa/gwC1THDbprZLE/QEvqDyTtK9qANayLDldoBsHgqnPa3CnZR8cSMq7p2Bth/ohiPfcOEgIIKJ
+YWoUeTso9qOKwnO0l6JOcH1+J6KJWuFRhVvb18RzTpwuFmSMPwG00k8iM3wbpEAqZrglrfisKTd
XiVe6xHa6wgF4xroLiK4qCQ0ikr8eAG6KWh9yVHoYTRVFHXAXXVZHDkAa2VVEUQnaJnaPG8jnbXU
o2PV8RhrT4/hfVsDGTmrp4elNsD9O2So8iOGqa9VYfHbKjqLFYTJS93UjpppzAD+XLJFh11AVDHd
zI/JFd5TeYDCrRufGJd9KTaENZtJpQaavCovLJHYMx79wJqFFEa4fRg14IDpk2DVn+Kdm2iqHoi9
/iBNb0hjVKHOy9J3bdXouRVRu6jUyyGDb10yRQ7eNDf0fays3KEIYqlD8wKDeVpvNSgiu/MPBTH6
H8lZAtVUr0dcqHtR/DlyeAODXj7GaKycNgDZvRP3ue7X2iB1GDpAsVqf4aNm8uZFW9G1/uZHW7ET
FyQX588gzSA77NHfUNI/5VWPoLrwYteIHPTpLkPtcgX9JBU6u9AyX8JS+r5MyRX8DmmiWWYqm8Vk
BkcvAY+0F/T4rhrUTv0GSTRzYfC8K2kwK8JlToIhSY5pfLNlGzmHHoCDfkubRsqCtx/7Gc9F7tlk
aFN4I7BJKuRu83o6wslshvMcbRdcgVW9O/20ZEOj2dWmMieKlbIVbQWuf0kTmaYXbzoQMYi28uYo
/i5DhhNJmXDL2Ndeoqew2yq64wF2/fcHH2DJNK22f6KcY1i0eWkXgfwujLPNx2kZMj2d1+nHD+au
qTb6zu+OMdbzUyZFHGtwYb/B4gkYWwxuZpOz0ZcCR2zZv5GzKdrC4vaflw6C096nvHEyYP3Zy+xt
5HnmYidWvNX5jNCydZs06N+w3j1RayJ1xwji8rT5YKe4UmWPFl/dQWEvMYh7vpv1y98+yAUPwSpA
LerMA4X63WlnfVgsyT5Ro6+AjB9Ce/3QuslX9+SlVs0OT/z5kxOcIX2v+lIQvsZZ3VI4rvk61etR
asQTGr76JRhBnbT7s3pOhVq0jXDNnFFdbQjwf4EGg5cGMBhKmHBFm1FfD3hnXrs5A77ptLhaPRMc
B+07AedIVTDnfqhKbeDvTVSzbByjPlwjeuDaNGzgcDYHdVAQbDI6rnptV2ZDVGFs2rM60VLvBwyG
YbQpfiBMcjlIDI9qSmxJq+1qZk6QtmVbj6CthHOKdeA9MXaJVdzPljm0rgVADS2qZlkN921seS2o
BJ+vdxJ11wH6p+Pt6J8bsZRp4izswV9nfdI5NJ5s7qDAAva5Ms/f6hSBSjX05SsLtlyPpDEytDCv
em49X0XgxKvqZyzQO7glCkFruvTqj1a5a8BahpuPkYfQjUXqSaHRs3feYWnXJtr2jm3VV12a8oBc
5PCfIZslKArYeys8yZ8DtdzellMMY8+5dDKyJOpar0Kua5imSf9KtWT/kSIa+2JXFAPms2jQSX5f
4FZbKoseIDAmNtJWwmOiN3wUcElaBssIC+v4wqadMoq4FSeawgPustLyXSL0GlSjFBKeQCJy3+fn
GiDpLv0TcrkUlYxShjzgDuPo01gAKZewhFgm2l71qljiy6GmFgS1eVzHhnNjpNx3GgIVR9jVHWug
uRaJuZmokX/kAeg94HvupqCZy+gzKaLhQz9fFVkiK/r6wRAbGGUC2wQdn6qPWvJSZFwuiw0lBhoQ
VfBO8+PRTBvlxOmjrMxWjWRFVSRcm4ukT9TXkHFUfDlOFiEqZ3xHPydraOAVhl75N2fU5L7d6jg8
6RCSQGcVYa1fw1bdfxyKUm8AMEoVxvq5bUsKPQw2Zij41t5Zscu6nfMED14xUU/4ZmjOHEToEgln
pA3Kny4s9NuWkKJlkp82f6eN2Zx7w07qIky9G5/Wq8KqGRedoiD97PPUw55HhpQAGrDQHykujuYd
mQ7R1pZEezaTzLXt1fBZqwpYk6ByhLwfaR8ur4L82h31XDalscU1p6SomSADUvr/XTA5ifpY3XKd
VpyB4iRjSmpFspL1AXYIZA1CE+rZESZVOqUyhhWeEY3J0li8nKlmsLCw33fPxLFL/9XhViJlIjZ/
tEwXqwgFLaz+6TAu7J9XwNcmQjZzxE2YCEkeG6tBLkp4i/izlNRlVNiAdjwjmUM65SzK7Ox1fBBj
8V9AbucH/HChvAdJ/7nIqZUDFfPjG4UmpmeScK5aeFuz399OM4PM7iV2KBUlt7GGJOA8+08Ph/nL
QUiZWJ5ln8+eLN2KQYCX80wm9wdygIRnwi4ejul/Q0+uHIam9jdwee1Exn/23i8hkq7Ff1YBX1q8
TGC791cNSJ9yYtc6iYiN9DkKAn7pk4l9KC03hoWYJ5IVn3OOf8SyQ+Gf1bRY8ehFKchAPtj9ln8/
E5dyGYkr9McAC6guY1haVbdTk0yV1PEE5D8Jp+XiAkXrR30KyieWQHrwFR0ouBpc/vOo2meUAa/A
3fp0PaqOA2JQXsopYUCj1RnQovlqf8JYOGnjBxgFhGaGBQatX0HXRW0WuNx2z4e6qtATkHh5hYb0
p1jBJ1Pecl1pUBWy2GsOzLV8wFSGGejKnY7F6NfhD7NsvzjXqWGNuOXIQToqbdFQjL6WWLahUBtr
c0nW1vNF29N12XBJL7H+Mo/XU2PFbOdCHJaxe3paUFP1lqmBGH5D/uKKKFa+ntV/5ffoWiPvexDh
9jGcUn+2gYn1Mv/IcHYdO6xySDBrWxV6IenC8aT+pSxwS2PyaAHTi9n/+T2SgeHYc1kBWsqfU/me
SxGD2lXH1/HDNK3waLHFJkrvGwsNK9LWRya3Mujye+muOIN+cUfrX3fis+vn8GPNgWvWTFfcqQxy
Fd3MI3vatI/VploOZbwlZBgLGdh5RadRw5v1E3I9vGTdZOVEEP/wEqj79N/XPfvG7DffSY8fQT7V
vWtao6zWDoEFCx0uU7lte5tx6cltRHhn+BJkVAngWY9nYfEznJJJa+o0mc0KeTGkQsVDvIzAdkHO
4+nEMMyyvOQ2sMcA8uP6/KqW8myWi1d/qNLjRWjovlqyLNhWgEG+NArkO71hHaNo1X7maxe5JwMY
IrXIFFmldgyrYXP0QymPjluEq+heSmgEbo0B25zZmqhRtJocRLWeAexTnGg/SuvCtk5cEiaGVNnv
pTbl6pDq2uokoh6xmqoMGlrGp5HaKUgTW/bIlF9KnEtq9wVMKuJuayoYNmKQNXA17fJCtJChm23G
eGnuocVHQSuM7Hv8KKJ1U0RiYOywAhtfOTXDIITnl6lzrT26/aHlshecmG6WLi9wUhCynCLhhfqY
ii7pAOo7yuefFAuS3nNNH3UEQyJzQu9DJit75UCO6zU3JELlDCZSwEO4V5yMuG2Ts42y5yCVuvje
Bb4QGBG4OmXp781P+5+6/vGjr0s1wCw5kFTyqC/bGmBZ0Sho8q2ER/5BNinDahmTXNRVc+W4db18
nNanRMx2Cyjuplml05OMDvOnmj+wXrcIkdrDPBWY1iaipEcu47VLvXKNDr8Susos+mI9iTBqOzeW
tZcvPCXre2+jXIi8HhCVITV3hdcXtVRs4kjxJbrxJ4ZKQEtZjDsEqfwq+vXpIuFWwUOr2vdhWyXC
L6ya2sw8bgmiVgeXeL7Fj2PY2PYz6xVDf8J1eN7JwnJUSyqn4Rnmb0FzuLs4rj9NjR/mC0cGnCro
oVchdm2l5k8TflqzxfyERga+ietbmdZ2aYJ3fQOlhjhlifSHAOzaWXBb4/WCBxmloxGn9f05AP3v
70OmTqw1i3kjBncQ1aCnrmUAPzQ0+6z27v+VA6LLmsPAu3hJZtD46QXHbdgAmmnCwhMSvZhpVtMT
x7aEDUhuTphFnxkGYQzEKm80NfLgWC/wOOPmQ/j/cWfgQop6tEZ770LUpT0zYeK2mX5nh/jmA4Zi
dA1/4DHv/teZq4P2WIcZVAcaebdL6eDVLKNy5T/0WXSgj+u12ehxFmwnLIKHAiRyR70GRqq4vwFN
HAU1R1OIRHK8a3hzG5vk9rxI4wLfcjr/txNJCU3LuW8Lv1OWIPYM1XbJESUCECwwJ1KjN4tgo1IN
nNw/xo1vYSQFqGmYyOpMX7L28nbi0TQSA1GZ5bvLGGqUZ8esH8c+BtepiHHbpM54ZhiLznZ68MVL
8jUG7Ips0mTln7vN/7BGByA7tsiXuEJedpD2SKXoX1JH+p71pzsn+dFR3k+pa9AmJVV+EJVc+BI9
VSzQq9PNRQSmmtC7TvPq8heLpyMk/YCUrNFG+2gz1xCXWrcZ9G1CcyOLclLpZupheXPxrWqb5ae6
UcA3CGN0nsKnkTUNlmDO43t9ey3JpEIRU3SX1uhtgO9AmkTccKyOm06yti3qOaHABPxX61FgMbvL
2jiQvUfR8eorc6zCplcI0lX+Bxf7/fRgkNbnhIDTZhNnXeA1ZJ79Yai99MQVJ2USwQFR3ShpVSYv
8qutGU3Gbz8YJU1eK+1ss6hIL+BlS8EwOHHYRVoP/WH/yuInj7bwapKOWKPjf/CHybxuBFlUySgd
MsEXhc7wBoQVzqo41nL1mMju5D1P06BvTL2r1fvVvhMZOJW5+L3ExFhN+c7YsLOZqbpnwyioj4gK
Bb8xZAvGslCkRoydiR+rKX/axiSfOpiTUsnQpSd1F7G3TePrEkYuBCQcp+Odh0F1gsn4wS80IDCz
Qrf6jQp5bju+nfNlAvGJp8BoOaVdtxXdchoyZxAtSBvNcFIP57946rEKrAcGWpSuCyCGTV+FtgU4
/OUfv+NcIV5SmzXEyuQVgqIisQm0mBOCVW5f6RVe6mtur3nSYczon3HQJtQsUt3vK1jbaMaQKHnM
dssgEwlgIRLhQ3FIa92E2Knz1Uks86E8hjQAtftb3sg3+qKJXDfYsXPumTbxv+K2j7nARr084Dhf
Cnzdr68rUAr77tjbzNtVJFD6kQfJuwRH3oNncR1p87U5HT3XzikNT33JJmePr+FKPNaDr7kx0B09
dPjSkUmhDaY/Yo8tWdskuMHgZ9IcJjWbFMlOXxIxg/J8/6Wzp5xKWoZPnrQbhBDtoXZAydh91Ogm
ebo92KCM2QpAdGZ5tsZEj/sSWnM9FJXCl1i9jtgnGcJTUxVAycPrdXIKw0oIByzs7a3o1Xepvk+a
v6j2+pKxhuEt8+goFq/eipsCuczHIq7p7fC17IKPxC4obV67r6Lt+HfZfG6salchmzwtXQ/BJCYy
YzO8X3QXRdFV3QGb1faZvGns8xo2E2rBdjluoY0FgIyVKQ3tg3kC9KlYZb+TKz8IxTrdSzmcgpCm
2/uN18VHqyvQwj0I2w74S6+E13zYn7JaigYJh7+hs8JDAwGkcL2nC94tC7skKRZtIkbZx8zQpRsv
IhsQJpER9NoqzrikO/DU6/eDuqfd3Fdb7uQloToqzQ3VrOsjdUcUyF8gBt7wj7fOdUYc15jjvAFm
yk8F9ndgXbJfHzgHpXRRiZuDTyXQ5WmoT8PfIUBM9FLfhZabAohxZWgKqwvCOh1ZNUy68nNYhTk1
QVlNOiHA8i5NKtCVdeIW0+j8P8X1P0rfH/BYgDkUeQVDh84X3y2uLdyCzq4XiWf41iO8JEIRhiys
trb6rlEr/y5IuCZou7mdpKw07cfRcO+YyGh/zEHS9FEF8e0vk9mYVNXzPLa05fGQa/eARanjW/Bx
idS93M+v6RozeyBBRVOoW3ziLr40OXd72OBoYBXD3JWVr5EJYcLgmAZzjk6H41Q8Y7XYfwd57UHp
MZCR4lPQat8LrL8FralAamWJ+6H0tMiuKZRxPavifqGyTfJRb/PzA1RydYWUHJzewla4VA6UoHSL
OkKowlq2warfqjN9sELLj9FamYsCI5fx2W50NiRqPonDlszEfyn4yrQDaj/bchODqlZzf3uh4YnH
hoZE19CKnwCxW+PQguxdaJ45vTsPrGgJUKSN/gvGrpil0HEUv7zhjDbe/mKHthKKtkE20NVVAblI
2DG26aOzaMpLVUOy3D+uejZGHnstD2hzQdYf31zpDH3VJHwVSBDGPMMp4DG4nP7KBesb1CibIqgj
8PalJLvmHeRV/Q28FC4CD6+8StORyxTz2rEOoBAA2Y0+KmIiiAI71keR+o4Twd0lN1m2ALqOtuFz
A6oUCI8P95dRgey1LEPgG0qB09XaSTop0H/NeyJWaX7zvibvKfP9e/+Rm+vc+xEQAceZ2fR5VT7h
USMZlxQs1DjKJ7PrxR+uHhPLHUvzMUsKqi20y+45sy4Cf5xeoLeMoRDawrBpfcYxQv0RWyY1KSPU
XRfxgqdEU0QVGeEGB73v8Pl9hv5LS0ZL3hsDYrRVgaxJ1UGpaek9Y9JbZ4LuBHrS9d0t//wfAD14
1UpVd534zBxo+XxRRk2+qJXTg9g57YeyUzH7lNA+95+tRjj22619SlytwD6Eh1GU+EDTWqqCrzje
WbaPKg1FCU+UTJxKPrDBXknGLvihg4qBKlJln+FVgliBEHm0xN23nWGWo+djKvfaGPFu0zXtY6iv
e1Efwo55fpDHaNq8b0HJ7fOK4qdl/RRBeyn2XtUGnuf8EsW6dNPKyEUkLUUJfqqNUAsgfPUoAKt1
Ue9w6ZypUv5cDqHZFjbGWAzwBQX2zKa/SpjBRGmRJs/4be6wSWXK5OmGRApOuaCe9/srXA/ipcp6
iYwAtP4Y3eS0zaLh3b+3bxXxIsCoZWMGOKtX5qljz40ftys1eQ/NQBgIjZcEAeS59NobRSARtgbZ
i/RlkIw9Lwkh5LhRhNvyqzLBoYLatgGsGZS8ytfuj+K0rEear06pjBTKEJ1/xybcRaL865Cgk6oq
NsY5TQXARQC7m1f+JjqGXd6wmarH68ZhLLq1uSJlDEl7BzpxJGmgxcgmiunnAZIzWIBNmCRYDZtm
qr1xXe7KnIlO+WLPr4tsNKHG0fGme6jf+nyyFHsALlq1/ZIalvvZvtHL2Lt5xlq1DQwipZyjB+5i
mMftbL3zj8KqHcotrg6lPTyoRaXsyxyJ5LTeL7+8mNdJnHzmkw78uf3HvjoMGQT1XmVxEv0+5BCj
sNOiqIDMPjB51AO2XmvaQ/I6OygQ3P3/fdNG7JztkTNPsGBmrPkqTVIXUv+JO+guNgmmjXdnoFhp
i+BqC42YIZQf8O7+dvZhbvu9DB0fueP6T7I96BHorJRGxMp+TXUFIqgkgC5aikZTqxorG8IyROfc
yDOWr79VfaX1mb71OBA1ep0j6pMphGIG4tKtUXTwszIJdtdFIM22q0rM/fmPTEG4K3QVDN5wDzS/
gC0bIJkuMG5VLkB7LRgyYlEPhAiwVWWMv+57zaYomvR7Vb+4nwBmTpe1AesNL+Ysl89ZdSQPMgOv
9taS6GTZnIZvRv5zRrfySpemIlKsKRWklzwk2zjAFZnXw5+XTijt+7ejNniEkyK3IPZi562Pnp4m
W1FDFVbADdxPDZDwgNPDdlyGKD9XXiB4zEqlB7x1oaHXVyOVx95FNaQIFU6yvQpwbIcvJ5ObL50H
jU8mTzA/6mT/c453zFeUAyA7ppLoVUy8GZ+3WghMGjtCcHDfbpLhI51tNFGn0NIKPUjQwJeDSKew
3fjnO2BwHgBmKKyzv/eIf/JvL06AzJIf/q59X01pJ07LhII4OmVKXlQrnxhFpOnEWBqHsjoijWdu
GHpwSXZjzfTg+RpPrBLFciQX9UuXBG7aEY7eEbSYCyebizOi+bf5tQoLxLJSI0nTKIKXT1a5ojLv
wete/iYRt23SajuDB0oYd0pkLjlQztpBzT+3qQVVXJdqbbW4/pXTctri9J8cQU+S3NzrdSKNlZN3
lhv/Y24Lxw6jf/RCjMSSCCK9+D9Okc0D42s5U5KHs3deUiKbeb95ZTdRURcKoDF1A2VFDWfzPFSY
lbijUEkpUXnaoBrRAeIr4Gey/50XRZdJ1uoLvWDMnXsGpqmJXGg75Lw/e+YXAKakCSUYWXhgV8nc
cjA3gh6Gled7t0x6drEwlZhyN+de+Z4sXf6Mw3Vc6Y5E/4g8cbiFGAvortS6zJFFOSOvMG3f13uI
NavCuIy8ea+Tlu9If/HIbldjqwBgpoS3bJAaNds65MAQ574hUERVre369G+yQVajDvUKAGFUd9bu
au3yo1uEWJ51xs3r1ZJZ9Gp8iPMegR1+9eO7ErAv7djjEipn96lha19CCItAsQudLa4s8XPKoo3k
INIkGHzO3on0idy3VeewqHk57w0WbODtkbgjrNqtXhRo4HItMlWviv05y6CK1Y2hUpmVebANqIiU
bQ96HQFlzw7m27JilHuG88q0y47OjYLPmZmLzhmH8VfiMa4fxquwFrc9J4aC88QbVS8cot2o3aoZ
oXyNWAuQSxwzavtouF+LxsVPNmYJVRY67DW00F3/5vwN3GhlWodC7OdK6eS8HGWwtxLCDrkv6s87
SamCorDQApwtMuJLF761gUQliAgz5jeJbIyzn6qbN57cuyCiWkV3TRlq2fTJQkWPNR6BYKg7W8S2
pylcUjZnZr8ab7RXefDCwMqClFPxZoSZsAJHjZu7NksDJ3ONUeYwKTlZ7dR2swe5ktGNDmNENtjK
r64i9M1N40ytG2a8PV7hbkJSxIrUkjlPRVbs+1sTy4RLMoHA97GLqSnBkvUyFLOC9MWJ3tNN6oLH
il0v1UGyHg1TEM98viHqo+jIemLCoMWUiSw8RuZBm0drOQo2Wwcug1kDCZVS8oZc48SFHbO1h081
aNLZXAHRAlmBJ8c36tWs9RShTy+kScCV8Qrh2kS0UQIAsT7iDNwiKYMmhp0uxM/w2RStc33k2MTu
lbRworCpmWj9J2+HaAPeqXEIfAZjCmoujIvzXGtcfB9xJ45W8GzPjSTxIiiOgFfQacwt9VVifFm5
6iecCLuU/6l0+u1JF2EDJtIzQNf9aM3ceslDjzMJo9/aVcS6G8YZ51cxYOyOorSAyTXTPhvutlhR
M5dFNDTzmIzK9RD7q7eue95I3KTkJinPODxFyJPJYl3cMi7UsRJLEKIGW5q96hwGyHOpAkVhvLbG
DGnRkS8zwfA+qHwphA1UWNIt9K7IIVxCAs+I4WDFD8qqTXbn+vNOymlYrDvma59Y0CC5TzNbjym5
fmwX0/8Ngywr5115QSMognbcbWJTskLuenzzMwFZkG5Nw0JDPFOg4i32SPJTiAZLNGppg2bjO6D8
JjRz/jmRGIcFqif5U541U6K5PrO7v6hY0OjguWU75RBZs+96o4avhrrf9s30fxFe6nAJIOqz5VJI
IVFY0+CGeVK3Xz88bKYq2hGIlIMsW0D5X6w5ZZ8DKStMKD2speSTBq3nNfkVxERCfteVA/zUCkN/
wcUH3ENM79sGHE5q7krW5lwdl2Z85l4xF8X7UEbau6rYFWQyHRHQa9EJAU3Jo1PineU7IFDCTNzZ
s9TB8F6I74JP4ytN6YQX92bJ2M9KMzWF4wJBRpIj66pTBQxC+pYSZih+/MkJ9Q9Qcu+VW/7xIES9
kfDv9AFKviDa6p1ytDq8leTJHddI/ZQUZwGPRuMmTLAwP1ObPrxjXnG6txlNJydMTPw6dhyNbEPS
LnrcGNCdOU1zq6LCpSRMvhf66XNyOL+1z9hNpvIyEShcfOgvn6CrA0z2mGvc8qF5NA4WFd06Xi4E
JnqwamyJBRlhfdQfTLjyaPFx/uKCn9TF0pu9Y4TWF4LMSwVG2AyOOarKcjJf5gdQK6ae5v3QIGJU
ZLb0fPOh1T2OorYkzPCkm+4LIwFmaPVhfIUR4ad9jLn4mc55cB1DT0QSdt7Y1q3NR+fMpAvw630D
sIfPZwVboiB2zBdYvPGhZC4SaoYNI5M9Ly5+MqLG0mmm4CvBf/6vyvD9iN9Cv0VmCKJcFL/badtT
qNSLQm3esaDTaLC9eAbIkqPrvDLKO6hnCVA++VKKTeek4pJozsz5uLIGQ8tddh7P3psBbloR/03n
wZ8sK0XFDaMhitGQnTd1mu3fYgVYI+wFiDEVTIWHpwxBbK25SLK3mGV2RYHfeYH9G+ZVhGyJS4YX
poRXMxxLgXRghKNZ2Bt4YqfBngl3x1bV26creiQR904dfuvJ2O7WKHSGQ8XZdfxMYPAktb1U1q0a
vfof0g1wo5Ggkd1kV919YwS6hW7B3VyhhJ943t3poR3W7Uavssm1rA0MJAAhoHQhUEzPrcaGY0mJ
T/IA7/E+ibO6Tmzz7DpS1YNZpxJzFgixH5ZCkEaJS0LtUSKDNEKxUYvfOBTtVhmAR00nJgI0et7o
/LP0Fnxf0KgH6mWWgZmFGrACjTkaVTSTNj/ind4n82RZ/xUP1AfDCdRvXBLLvqkYVceusmpDoGPs
cAN8cm8kIBGsoxI6T83xQrhfgIVVxON64D/cse6qNXNC6icFCuDzgtYZjmq5FCYvUG+MBt0XTO4B
2CTIyJjhDoRVkVoTQjRPCnQm01w6jZdpa/CXB/s6jP15GtmeLH5Kt5Q94If24LYLD5dHjUBLN7Rd
k962NTmor1OhLaW8UubVWSdsoK42ONRUbWMvQXd9Qem2y13lVb9/4+N17kGZZ6qHahXA3u7xfkwx
W3kkRmMGeJ38cRqjNQMEcu70JKf8b+5lsILs9q+vvkIaNrTlQeWI+0WMsdoVEYda1ojxeZUB1LRm
Uh+QNi0ur12k+S9aShHDqH48Rsk0fNq2Qz9s5TpVa2YECCqeJZo3+0FqHNd+7e3+d9cgS9D+KiI4
f88GoVbCUc/StaAuofPGtNwkECeawpUMBqUWfjt5Er9FJmf2ZQ9IOU0ffiI8sxJV1uBMG4bfvREV
ttxtJtaP+sFTl3jxVl8nxQz8kI4CWFVgP8QUjV/ZGjizeH9UtrLpyDj4V+BMtb+nf/E2ZaKpy2Zl
lo6CclF0oZG4lkNG5DXAjSzr/Txar+HBr88thF0ZElkEBdiN5DUAq/iyteaOm22zp6qWcsOyNsCI
xULPcK12Z07I1vN/971gN7Lv3GmpBD5AZ6UYiTt+Ni9otGMsZUWNzXg4vdQXgNbQl8TMvsU21F2k
y0+tLPTmVgJ9flERqmJy5wppjQCi5hzWwgD/lI+AzrddWmINYtfVxsXjB3zGl3vFrYTWmMhgTIi3
yKstpadzZcKM/guWW9R4pyW9DzypGbADp1ocKU7++mfYyE108yD1wvxHrOMXryiYu4mmAUkKs0sM
qbiQQyQntLNbK+Mb+Zbjq4L/ObghUfTJNNDJJ26wYNA2P33oQmaAJo5+x858Av8kBdVVjN/edgwz
wuCla3WsJjFOVm99bFAhxdIq8rrgWmWMtjhV81rxR3MngUmXBIuBjtVVvv/PxAUEq8Ipceq6twtq
7EdmNyIf4JDuQ0Ci9A9RM4L2goPZncdGOoBiFhMJq8GcCrh5cg0vn4xmPJ4CRAknvRdrSqT0DuEc
cLEI80hjeAfKmgatWWbLmRsL7i6D4VBB6zZPn2qkonRuferr0mCI/PlaFSOo2qrOnVhX+k/nrrPH
vpF7a9CSzmP/qXbgCzcmJ504F1b3+XcF1aUjFyE67EeC+8Ickp0bI473dFeO1+tOvOxFVHUC67hZ
HYZbRjAyotehYdwyPoG1NLn0SuZ95nBgJYcLufJ3GoOslSiTSl0DhBHB2aaGjligi++ImzYLYp2Z
I/fOJwwF4jPbzb2Dju7yMaX88itMevXWI0D/myRWuuz6lv/WnWFgUbVntWERLQnSRH73KOfsSJ+v
aw6pNdcu9tolCcqO30Na64iHc2niu6nB9HKzWDxJzOlW831fQ716HcZn/D4qukHTw9ZAD8n3DbMf
EGD6Nb3i2UmXD1PD9f665YuQyD163b/8yrEp3Ve/YhhBzs48rayyZfQ9AIiMh/4YzhS/cU0hyK3V
/C0wOZ9oi6XaFg4jDLN2M2JKWLt4AFKC1y8l9FzEoQE1+onDgLGO3tA7C1sM/YfG+g50thcP+qnP
dNK88YpL+8rUzRNUNVqZ6xitNG+Eno1hxzMpR/U4AN+Pca34TNrDz6kqW7dBWJn3Hge5vcJuaCP2
Pvu578EPYMzio7bhsrXqLjCUQRn/S0VIoHbVtH1Sag8FuCR0Xs3ulzPvT+kJ8Na2cbDcavCul4W3
8n8QBIYdVsmLSVL+JiNnKI3N83TEesE3VonzUZVAD4nNLB/ZG3ln/OHr7eIQoe4HKEvUVpt7y4T7
knmwx+JSA+Yu5j59JMgNKVQ1hHVS+xheFiLBKJ1V8cEA4EiuNSjdnnzRdBcGAgyivxBJK1RmRhOT
PAz/mJOo4EliYdd/lSeekNfhyB6FvLxpQbEGIowu5PA8vMBVL2jKNYR00yNjRlj1pQsVS8GlUxHf
O/AfHALN93OARP+cN2BHB+p1QcBVxWHjaAE9zYLPDnJwEUY61Q7nfXmxpkMtiF0HQpLZthFlioL6
p1Qd5+HGOkT2U4lZYVRj8RSWNVrQvHgc6O5Cxgny878t21OoxZSqKEK27s1jyFC875XujWEMmYUv
kJGR5vIUEHxFedjauxjEaGkCdHOdt/cll7K5mvUP1HTjf83tW8A/V34AVOGa+9T97tHE7thgnxn0
PkxVmgKNH/utSLLADtNzLM3kAg1lV6B/SKZfBtsNuHGglTDcod0bOC0lxf10UBsxnSOZEkdPjsPD
hUDaR7DZMd3JDY2wtA6JOLv2RMaYa17ec0SGseHKWcrPmPRNzNZA/IdNDxENl/og+4Kwv87fBgZS
yNLb+kxEdf9/qi2ILMfaFGlx4qttvmFlLRi/2X0sMHdiyDHnuL9X2KOIbZlh9haFPlQ0IWgvykDk
cbiCMHr8IDZ03ZArjuZYSGYH0OFF8j1CT8iH61TQ0xHGYMEnMghaqc9ECWMaUChWHj56xSR90XuE
Plhc1+KQF/78jDOsZbBPYkSRyskS0bN3dG4n+B+ku3t+llPT9jsqEDIhwoO1hbNbEeUBbqA3pZC4
2Yj4m3yUpehBPaDbFrKcLltnfdx6m/OrkqFeeU/nHirit2E3nFjAGP8MwnMVXiXzySh6zor9yXsu
A20Z6pN7Es/Gl2Ia2dunwkYQw1sqPBrS7aPrnHeDKsWCQj5sotIeGtz5TCJjAS52B03ZsxFLEi2J
C8kxEYdcWdXF/WRtZvFW1YXO69yycMrqkZ4/i96BTCBSIDnaY4ajzWr0klKcIRb2SYyrsqSfabEU
pHUqYOTs7sxo4TQBUG7b9vvRjx7ZDxCD6rLcVUV8c1bz400DMLthO2yjwL+NlXu2rOxFIFLeOfum
Ddc+kUiUNXdOuN+jrG4QJVNti6vytDSzYApbqXi+k//h79cXkcidJ6e/XeLqkWWZTlaVQi5Rr4QH
pcIdcM9gBxxfDs9rSo8E6cQTT2lfuOH0jis7NgSKxj/Nhe2WMB4YeF5dsGHRlRjTbarHpcqUg2Ew
xZnl/N9/tKychSxJLrM+2MFJQDHvIyo5pDYD3aY/ZLQMaaM3zxCFH57bB2r5EjQWeABMWkrAFSc8
wD9GQvs9Fg+qw6Q/5yT69K2xNzGIkQsMSmnGz6wTWzMxRwKQi/gDoqIbTy3nhTE79jNTtFUOR1tQ
G9ubnHhQjFQeb8JPO3jUUAzbLaQxNkvlq0zdM7/fAcw6wuFaS8ZZgvBu8lhKuVCVEKVYcG/nV+q1
WlmkRFOWr75ITlLNUYDH4GyH2kt+YPXoA9ugbNxrK0FD0GBvuMk8h44PcjTnNVi9BiUX5RJSozmn
gZrCSot4FSAcc/GegqSRxE2dsPQAGHMA0LxCKBtcsH0C6Xrv1mLNeHU8LCMgRrla9bBCRPa4+w7n
bd5SzJ50tHrsgUug1bAu9BecSItiRLML0Sg61yh3QIefYpjptPjLScO94oRT6F7+xoP3kbVHrwI4
qI8VdO7IdG8Rlj+BNenKhZEhZ1TqpMOW7n1OpwqsQGszLkOijSSDQkrT/NqQK1L8t8WgfvcPPDuz
NY9gUsh/VXyt7Rtgct8NMc+RiqG1wFmmqpj6c5EWIornNGPxfJsvht++GMBkke3dti7MTuvZxr2E
7jUqSprgNuBBlIE1nAuII6cwMfyNROoZ9ovYR2zg20/V7FyrxswWeAAlppcyCO9ImwfXXKjCMRtv
CJueQoVxypgmlGrZbvzC2Adt7glEvNVuyjmzsetsZfAZ03+9ThYIWFf77bueGbP/OISrUjpCEQBM
hHHjB6g3JlT/8QX95O1Um1JSa43J25cZ0IsfY9SQ42qZBI5GDNJOWwyS/3P3wopq5krSZ86JS6BD
GUsVsDIk7MpkW2unpOIGBqszrVf7WzALabGomZowPvjc0dQ0c30+S1QXE9lApxY9JPs+lAIxOolk
ApWyAngKDlCasm90VS3n/jeq+ypUzF5C1mZT8uhKKVZCTIlkpMggs+AfcuzC2Kkpwu/6lY0EVHxa
lPC/PHZOzmuw44ZJL4LWcoayMuLIVFKOJY+l8NXMukhSHlBiUINUkINXiAKLsBTkhSZ3PoEUC3wy
ey3ijjGrVMxYjLvO4j/n/N7YP32d0RVdX423fStKzCrkqFhUOY/Z+vO7EpiqSwwdhV4yAH8u55z6
fJHEgF16sWu8iXTPWMLnhLM627lwiU3UOepnrkkBUtKnvUNxzwTQRhD/6N90by3+LONdnDkXeeGt
A2hOAN2KqSKtzQYmpQayhlESCZjbMiJMtnlRDnHqv1rox3t6FR9E/1W0TtzxByQTfjnzzhduRIkj
nmilNmZ5aWEiUEzWkwThUpOC9IGlzjRPiLyISbdnhkxEQw4pkHAYvRM5Um+vZl+DB/OFMZpxm1Sf
B9xyup9Pk4q6ScQRcEkw46q/lEVe1p0CF9aFPN4U/Ntc3XIxXOpuS6dfrpimf+8GKuKbFOYnXQ0k
SccAjcHb7F8j33jk4HViP5wtid0BhNd7aWJens7dkhpZZdqQgmVLIjaHjvSDzvTxoUkY3Qy9aOqc
Yk7RmDKqgrgl3XCaCC+PjZmLn3OgQpyd4NqrxMUrlRFFZB6IGX1vvS9b/AcY3QjGijOVkDgHGlsj
FjcbhqKAW3qlW7ItTMHt1xsbgpPb47NtSJxcoqrulxyHMO363hjY2SBv3EPGwSfNw6zXFm7GDEhX
xhxqUpiG0ITSy6+pnU2AW6Qmr5okzZGNv5JC5NXK+cs48rPFEl9uIkesLBNuBwvvHvhh//Jw092s
r76SPev+z97rprhvXwMI4NKDWq9sp7F0LYhQ5c2sokXlr/r2KGJWuQhU4h0g+Eu2W1tkLUpOVXRs
667LM4DpcX+4p0yqK2ixNT8E1RkheeITyeGRtqqYgDkdEDcrBCYBHYS6PtVZQjhPYHRRK6ejQsp2
lT9y9BL+RhUrym4nnW2NP8sGIWE6gzSGCouauabUieDU2hfPyoRbkRVQLzMSbOjljl1mKvF7l0eK
JcnR/PxAGM7n7jrAO/PFi0EK8A36f06ysc2XmDlKXfU7WjL6oWg8qb3TqZmH/91pOQ0ktXS7uSkv
bAuJXkdaIcqfQMainvrZS2VqxUNZLn3TTltdtp4u17+MWtpkrPQKt6OjSeqHstn7HjtMb6cDcUlN
jErlUgMlUNSJGSfjsoUsVvPwR2Zl5O9kLAbfrrnc6guwNkf46AGHBAlWnH+qn4jiRWvOgexm7DKa
ffLB5fAbZnUnIQaX5WY5Whx317q1GtVBXLEAdKAsp8ecB8/G5tJj5zvY13IrDNVMgZAAAyddqSJ2
zRPMne7d+KKDJ0Mr2pPucAsE62/5moq3eFrwIrHyQnVESfRyzmRdAYGeLltgqRUzKUCmBqPGtOU3
yp0bCl1tu04FuXbZHDX01xW8HTl9APzYHTYt2VCHgQg8jtVgp4o88GXclWWszjBZbQeTOGzt1Vl5
vWgspx1Q28UI/fKDFgHg77WDMKtxmyw0dS70RYp0eUZ82dpvViWycw0wBRQv9deL9bmbONQbw1Tn
fgi/BueQRraWWGZf57o6eNoX2qq/YXGwc6idTgwRhx4YhtkkmRONjU1dqr705D8B04tR4fih/huG
6QBI8HuVY4ZEYQpBPpZpa0Krtgoi4S0zMz4ufHBSJqVkMBBBqso080JtJjE0QPmaD7wEli2PCmDE
Ty6X4eMtHfiRZm9A8zV1mwIA/Y7ZmAEOgMYKbovGQ9161YJYrc5L2jEG2mgZhkaM21xV8JRYzFHA
0GRlbY9rAItRRJNlgrKuL5J4oskDVnqdr1eGpw7SIq00aIqLl1sSXUmYaSxE+a0iGQW3I8p4j9CE
kqjkWhsZcdJTRE0vwp7sNkLl8Yp/Ouw9VQ6ZGodEkqB1rJ2x8nsJaG9JYcZdsStOk7XtE0W3XOkK
Wnp+HNtXRjpP8U1NzHJ+VO87khmpKmkIpznXIK9QEfkIXeEUOIQtX3NjSBPKllkFhqdIngNLPJGD
GoN50qjyLGPU4MrOp5IJw4p3PoIW7bXYyiDUAXGFJd94JmnVhkCPAtsFd+KI3U7ETNjrDKb1FgVX
LhM2rWtQZW5Ffy4u6wEdGpFlumSpMSGFjcsvrssjYf9wh/kZWJkxTxrLiJ8D9RU6fV+Z8C0+Smd8
b9nBLXskqIcO67savZ+YKRTZvA78kfCB7E67886wADIrciik+CfuEI8L8sMuEz7IOxVqPnEpqXTV
LfXWfyQMW7oNRQ7qZvbwBzvsZ3YjbSA5vpFidaeAdtRD1txLHqLyLzwdlQoPFOz3GIytCXGQ4gNx
L/qOBMLEJUABTLzcs6ZD+VVr/+TVCS3PbJ+AEiei5sbYap/Z9o6w3Q7VMiZMGYv/18zADX0R8wNp
0yRrOn9JFRyleTvGTKUH0o12wppOw+Qhco4zZdETmsBTR5Z0SpkAD/16n8d4UJM3RoyLAZI/55m2
ZKU0Q0ypoVvD58ryUB1SlbwaWmvo3XnhCWIA4VMyXiGvwNv6kAwt62n0cYtBCwsi1N1a40r/eWyP
+GjV4na/rphtNE/ZvnPj2xbm1JMbcP1J/HdxRaL/M03ZkrIfjN58jo14eyZzdUZen47JvO8eGtKN
5o5XyGYE+FHZa6taPDIkGLR6IYG8WaJZXs+VE1skqORvIuM6UvRgjNAPiCFeO8L7kREDYsf9x8vD
aWHG39Q0USHjLrPa4EJeDK+HIU0RpKr9Mamz6Ihg+qpd9jXPYxvkoBgqOMk72H/vmjl2s3i9eK2d
InzjmEtRpJFcFOZJ5Mf6+0ZBloU7Adc1bZDCRiH4ih7MrBpqT+6TTp/Bj5xlbgVGG/ZtWsc3p5ZP
SD06zKtm5DLZZaRKGQ7VHDFfW+2PPzYLCpgb9KyzW1oQkezI4fk655QfRD7jedci4eb1sg21lLLS
uOl9V+Ii7nZ5WhGiyJo3nowsWE02YiOd+MkOOom6oRWAC+N7nj17ZY6+a6+WTJum9YWJ69msDYTz
nwnWET+/BFU8j0sSIVYMOrhohWcm6V1f1vOHFOsXmzUDvmTS+SyW9EJL3bZrFmH+VpSi3+ZiGIcu
+nZCDWzI+X94FK2I2lfeNwbKb6Y5RcXGGSgPoe9v3HmeARCxm6BK6dRy4Rm7LTvdlPzMhQS+GwRm
DfuFO1qjBJmtQBlkoS5YLGN69JvNktch8Tq3ZEilSSZr48S4zaPBFAtSnoUkPJpdc89LlHlqfTTd
y/xInHJ/fJpNiPAMfYSr5cFYecUOLTWtDIIkQ27Dc5FlzDfq403XkROHH7Nf4WNgxTP79s5r1Vjo
ExDaXaf6eCfvdCiQWZWp7Jk4zY9CKka6xxd9XkjNXboZI5I0J0WAJWMnkCilcdFwZlbMKPOq4tS3
8ymAlWWIBgWl71xMgFLg4CuGfQtM9GfcOmxSa0HIED7Ht/Gubn/1J9ZUthzThJzRc6wZGtlfjdp0
4qYITr40wPnKEQ9Z0w1FMRol9i/xKokIW0+lg3wgUYAU4NpDptRWcbGNL+2eMxjKp9jTSpl3Xb+X
cN/o4SdGuYzyQWZFDXFpIwYL/3O+KfNW8Y9+b7kMda3naFGzxIFwsI8NGCuwRTMhHs4YtG6LfCsS
F2D/EdoiB9nqAKc6bgNsB12xJLeVt2lxZJlOK4XApa78yofusPoQqXMOFsxtVHLxFVrtbvNGXQtv
y1ypbdUtmk79OULQ10P8j5aTE7n43NoU52Ej+9IyFgH+W2lPwUTQoUDCNYgiZL2s2QbOFv3eQzzv
M0SIvCc/DJtAlww5ofC5WHSU0QyW5KWJlFxfQqnXGYDut96UqdjmW0z6jCSVXC1l+cvAMQR+n7Ys
ow/CY2iEIzYLgn3+xDJ4/ZsV/1+ucffpfR7PU5WWyoW9gsGxhRxt6+wJnVRT34Os4I5YGf+Go+5d
IHIr0RQbdpODRdnFzsnFZUf5K2rtBKzVcmiVSEmJnhT2wa31kflIbzX5HG0HqlLFLX5LuZoBJL4U
Lr+gisVZMAVwrwKz2Fvuo/JnJtDChOEasd5G14IjD7YMEKXoxrnHUOxU9XwV1dOBjMLywAiBnE7X
feWtoSyImeWZXqIIPqsGX2JzOwiBYpFpXyC5KiRO/ydZeG6xs6l20CnHT1/yiYOs4WKiDrKJ0Nx1
Qs48tv5fLBysMz+EGGJr4WRkc7yiHP9PeJCGkMfJuWzgRWIgnRvPEa1Cwie2flixAKv1Tdnn7AHr
bxZHhUQGMJXsF4Ro1mA01W1UKNXUZFV0x3Nnv8c6DI5o9x9FrKu+a4AV8gT+PmfOivTPOv5ibaoP
51K8VHm4Q061RqBGd+ZLEnTZskwfSSEixkpcGuaA3e5n24mTa0NaH8dggTWOklVRkBIfVwEPPB6L
zmvKHg9UrjLkr0m7C2mCm/ty/XNR22MeLqiuiJDnc46xpT2lq57RJRDWV099V8tJ70U090sW5YIe
vwqA/3IgTpYLmRxVnLHbUaw0L0LWR2Ag+taB2hVc2S8pSRN25mFdf7Ofx2cd/ltU26g714p02IXC
P3jd0CzEGjFaKUxkV+VDp1H2hmXWKv20HD/wgUKWEw96SoAzX/+XYc+R804l1lbEEa5doIB7QvgU
GlzpeKsCDhXt38GyasN4lNZaSyxhWKzLSN0iSn0WkcISurId7R9qkZD+hTMNEOwWd50WopuT2PG7
ArKThx/3SIWzmH1iy2NPkU4YDolp57UaBppUcuLAC2lIiMP6Z2GHBUxDvHVzC+NZb4O/TYGe627I
DUTY9DeEoz73R7TDIWIk4zNyP301iI8Xa4gDQ8C2J5u9Ha06MNYPYFEolQUi7HLMiGTF3+QnCZ3v
IZ17ZWgofzr42psbdmiYwDWy5rswYIg41ZjagWxgvNtIHn09+ATbiRKU7aCYmvdlNtRPFLamdUfD
dP0Jr83pIGH8/0w2OpKiegM2yIjei4U1ki+MNP3GD7/CYu4tcfwDX96G2a4PYH40LCXffVifzue8
hhhrr2fFVR204TKfa/Awt3QL5YPXNAEEvrzy8uKMvKMzaFw7CX/8UApvFsfmOxfH8LMaTHqe827p
NN0z2KAAaTEpab4gQNW9ynuEmt8mqBtK6ox8ruOZPEKyy4wgB1PNxqisK3zuNR2z/iKJD4wgWqZN
wz5XoWeUBkQDQ0VP9lGVmMB1a4pd2ww04yS6hERzv+Pk1gVilI9jPyS3WQDpWi6z8iRTk23gPQqW
cehMZpACCEYPHLnka4QV18W4EtYLKuLfdgpr/WwxRBY2S1GGgs/8OWaJQU89mEx5gXLbQsSiQOiA
lZT2t4AxmA5WjjW6SkEKbB6n3DqcswwAUSWRYY7CwexxwbGCZ5r9+CzC5qlYSSSjjViTAXxBuOqe
1EIXTz1zsGvzaezDUFTPLXMvAu7SsUx6lZsIRRmfnRuFpZJnUjbnFzQsXtLsCD0/w8AdVipCzoYs
Y5nQOCslsOPJk54sVCbTC+bEKceNAoyH2h47hPJmEm4oT16E6F1jQOMK6vs/wfqrUz2tUtOIwodJ
QQ080xo1wa6CwCRGx/um+huTiKgFuK9hDTMTqMudtyknEx49pgX/0QnSkdGmy+VF1HwMZBW5lYq+
lGuo2UwJHLBLN6g5ecK4/TDHrVqr4pxHAow30OnnkJnrkVWY+w5oGhS2ybbMkAKQdomoVbBraOlk
DLMeZofRuG9O7MCsxfhIw9dW5vt/rI+qO2XVahPRzaDkvDSBCKpiQ0KCQS7TAUILMMKVZH4WjvKL
A4zXsoulnN6LS2bqVO7psKNMLrJ6LLt5XrT5Rxy4dq0w1XQEs+xXQSP0AcJhy0kNecVt0NekATeJ
i0VIHd7aZfwURFhf64pGTNcJxdmD9Ik7E9YI0jtB6kW7MDZ07x9HzqZy/Jf1zgNMeQvSn4NVgKrS
E7lHxJ3+5X3OXKM9DPCUI6u810gEcoc7e1oiWTC4XjKjr0XUusNmwGQ+AcfcBNN0+jaOoHdzHWVc
CUsgxVmnKINIVdFUijdKumrZGJvk7I4TILu0lCtkUZ/Am5UgMYDwjbiKEUcPhAYwIBAuQWvn2DNM
nha3P+MULkQEKToujAX3cLsfhTUEEeZOpvyytQnR5tdWRpDcEdfWQko969fVjYNOKIAW0HMtS7qu
2INbQoMru2A9y6HR5vWOy0DrK4IS6FBC0G4Zi1xd9zaZFISwnUJmF1ppVXAkIAP6qlYafphtq0Kw
0QsrSCwNIXdZN+Ecpvcd2d6SmAwivTEN750t7WA36DYFJSuMXLKuq9ty9MHM8wyL0g9DKn4Wro9a
c1/ncWxsrx/EdjmRDS78raFA5t1nuvrCowyjXnF+mjWTOcztqvfmDWC4EsFsF8DSvcCNOpi9qOFW
EsrP4usnZPssOV4cir4HE2VLxWwScUpHcbXre0OvI7aSwgZapOD8TwswNyT8YBI0DQv4T2rEOmey
j6pnNWLLavhsT85CBlOHbUumWcaq05UNPofTvsLB145WzaQWknX3QXlyRgOadUNOUHX1CaaqN3XP
t+Qilg1Lo9WI+rhWnJncvUpgDhaupE6ZlL6kHLWivaXj3AHKghcURTxZj/74NXMFsnAm6FNe0zr3
5Zizdo4xLrBL5jNGKwh5Dzgcl5aOYxNhxXpjmjN4OvK2zpONc0S+4ZKeqR5lO2tdeidRp96/IyOO
XV9jwaJZqiAyl8beT/DhMgGL07OoNCeeuuZgkxaXXaybPHVCebiLgcgYN3PxpqeuMWfY++ova+Tn
7LbU2nlCLmpgo1k0Gq+xLOp+x7cNvRYpM2XfPckqDSD7GDpD3ezfj8ikemqjaXN3r7czVtN3cquL
KJWWB/79g3GRXdVC4fy/Yq+7WS0UUMyn3paUBDWpYmp2bDuVjx1TgjfEeteoAu917b5KOlkxx/7G
jJAlvAGgHNxaPJJvu5OW9QdKsBclNpxkzKhB3EaCQ9cUlqyO7an2/uvAsEyahbKZ+1Gp7gq61SZy
8yRPFKwuVpx66B0/577E56MXt7h73oFDg1AWcVkSWXiKuhBqoogicYa/LDo+FjXWkSP3n5Jt8v1n
oVSHbgwTOoZrDix82DVELMkCnjeNvM2aLqA79V3lhfh4Z8HkEtj814iQYvYIMkmrRYHDIDhnzHrO
nbQ/Eudx3vs615k/g9WUQXAkoiOVEwnW9ZWm0Nms4xLNqae4DFHPMpfsXC4cTY7uDZe5ujdUgZWs
TRbx6dcz5re2ANrM3RRk6Gaa7kxFSpZ+MWpfTLGrQKsv77o0A4Vz2K9HL9qSXg7hxi3RcViTNJ9O
nAVM4Q7WLSfxbFRntfHUbeNIK0Ceu93qJ2/0QcEhuUdqQbWSc9chnMeQFLe7y0SvyVD0s1zVvq0v
y+PVmCWpGR0QCM1p3pAimrg5Zg2zGMJeJO5r5LJYV2Ys2nFfhm8UAQq+HpVMBMPT/xHjFW2nQNSX
t7EKNX3uw0uZ7uRid92dqXHVDXJdrlRJ26eT+CJJbGb3GbnNBi4ZhnKDf3sdUpt/YGzRnCTWYa+2
kDvoEbhdIBh/ERtAvFHPLsd+PiUXVvN9sejfMoqpEdgxu3jwA99VnrxzYgpXaOtJ6oJ4sZUuf2Fw
Z3rbhyu1yPZzllNLMDArkxEBMu5EWsV5OhTm/EDak0YDplwdX1nkSKBhwvCPWslXk6k2d6B01qvo
SMvzuoSqLLP1OMP4T/r+T31C+C+dxkYDFRSg+5773i89Q6dG0PUKbj5tA1pSm/jOjjHkwqiXvBbA
0SvkXQ/o9rpGwfCf/+YiUO7mSmNHbf/1UH3V6HDVW7duLEMsv+eekmsTQp8mcl3QH0Q6zl+Sn8gM
9/jexbhCD7SlUV7uLW8I+HhgrrHnCvcG+1/fH7ofcRCNd6CUcN8ZmDuMPauMqRK7O8cQ0ioRr8WY
WIFJXWl85KpvTlbplsyYS/qIegcDSShwtw8VSHaDrrBT5WDFtZyPeVAHlb9oQ8G0BEv/CMRrdxYY
gwPufOosGqipTFnJ1RtiiClpMLuUSTbGiJWxtr7IMaZ8x4qGwiniHXETe+vZj01kmK9U2nntsAxk
nxFW4Ndznn5/OOO6Wwz0SR4pdU4r67prMVlnRLJAwa5btf5Cp2Ct9/Mv5RgkOI946Wi5jjhDfI1E
uawCdTOTvWc7XxFEKYQlr/z3xQXsDn5qaTAUY+hhM716f9dnvkaFFeu5tc7A6FG28irI4bcDXbYN
EflrVdEMVgj1XJChdCev6a1JW/nuwHvJmakq4i3GaGqrVogenmmfjIy9VvtwVF0Q1uMDykpgzFA7
/8xp1w+XdwGVrtQFPvDHd79b2VUzoaZl5i79AuFCGY7ztMRhdpGrWMHEbB9vxf4VfbHDc9h4d8wn
CReR5s/7Yj1kfB3EZBHtzoUHSTzgxgjiQ3cPOzeRfGnTJ5nkcEz/kqyqvKONsTyLRQrV8wQHLzy3
My5xGS2dgT16wxU7dvw8cO05THbiotujrL7TN64+rD251c+xW0sxUGFOPwI6hVfM0J0fc+qwTGPQ
ayxxRPvqLBnuFI8x3QZB60/i3woeAUs4F8n5hQywvOaRKj84m/8uID4k5pE+Ye4pu4jq3qUZ+WEM
pF5GAHLO4cuVxuApGzY2kK5rZ8hZM0uyDUSUORjX63QH1ejBAp67OPBAzEfscV6l4l1SHITYk1DT
x/E15XM+DcIuVTkh7JA4NJrDrL0nO6JnYkeexKRGrmqJiH5U+QRraSf0v25OSn+fhwbiQODYbrF+
OW7s3hwKbWYTedjVQPwNBMVvFp6YvIcmsmB8h4WmuAKS3d0Uz3sAumUWc3MN1uo6VKioL18raaJV
yReVkG6pKTKeBgYh+TNr4wU2mIDSRFxlZLOQk7uxqVQNVDExoXrEIzgEGOPIoalFe+bQGWftHQao
hiH4OuBfyxIY1b/oRQcTQnf58eieJ7bWKRZDeuaOwY8RKMwnfrARU2BUe4gbieQwQAmqqQKZRzSe
R1NOhcu044N6lEOxc0bdbmwV8Epc21/dW35TNHLap9BSFZ2WlCWwcjX/XraB3BkEKPk4Ob9MKWh1
XijJa2NwB7m2RwTJOfYXpgmjS7P1sR0dA3PY3GTVvmyTe1G1eW1Fc3AZ4GjEfPD85mxmdjiji6NI
ImWOiwbXrMF0Eq8B3z2NkYGzmvebryo4TccIfQA1BqyxgLDKDNEz42+lxP/WESCvr4oOmziDNziE
4/NwKODPMk4bbMgmqT0IRuPaP9iaAQjhKcBGE5saPpQV8I+EAyhhaxBcO9luOhfZJdN2IAdSlU/r
9BNnlgqxFI2pgdIUySqzvuljhSAAdZi5hooM8fd5GwWqsOI+TV8434Mf7G1VC1csK3xJdCFSWpbi
ditTbzlnTpRPkGQNgolF36nhWt4nvc1RyovpjxJfknox95s08emNLQZjwCDWW2EWuSkY2EkmgBsP
WpOH/4DGouGAfS5YltEzaVLam7ktfsZh79oid91OlWnu6O37HHiqcRz7om2/cMfVw9g8dC/T9Jl8
PvKkOaljnSes/v0fnjxcaUPfjwGo0AQKbq/ODfoD6FCKaaB/47ORXD2LajcKbo8y/uKGCgYTmYMe
/rSi5G7p25qoUX38WARFnnrOmDHXNGglpuy57dGWNeQfYPK3DbCv02NIfLMPL1PHFX3hkD7K5mdM
ghgXorKVXw7k1KetKkRgplJ/alE1DQWQpXPxh1ALVam+FOvAjm6z49i07THjLil6Q6EQbSKCCIQr
I+zXtl0HfpbJODgr3fOfO/I+Gk6P9AI//G/Oza6V3ME6b70FimlT76HTuG8lB+na64I7aB5sJb8L
bkyy9BWfsxoMXlZBJJKgCBCzOqdHxMtQ6USSGZMyfB/oKqWFvBKBmvJq/yMuNREmgb7zGRC4AjWv
UuR6AuD8I2T53LR4+63Iqimwp0aKeuxB0nCR7EUheHCHaTqvBxQ1Hy7B9JsWpMf7vsmGlIGnlBwa
xTzYeiVA7lVVaKCnO67Cp4zN3MZnXchS5GtuNQVMBk3lbYwC6KSfcN3/3QpC5Tf/H8ZjdGcYs8EM
RjG+kpwypzXacJ4NoPhU929iXEUU1FnAJN1Mvwuc3CP6lO2J4vgmMDVBYVCfw7bnVxJn4z6KbAHk
Puu4RbGH4XZY2QmMfMmjEhyiL45EKW+qmbLFA2MrE0JpH9usuLV2ekP5uSOJIiq6J21zYszLuU8P
tYJFo4Vys5pStEEVYbXxyxUYF3Q1ytkZInz+cNuYLevRYeguiLe+XYcDzndQnX+3kmVojc64Cotg
WzYgzQhfZv0xA6TKYKcXeYhamsXDOR5TS/jWIsDVzUNdSVf038t3OmJmSSUp4cGkgW71lX4pa6ze
TdAQ2D2yajJ3TEW66I48/1W32XOcI5rKUIWwuHt7Q7YabeAh8XBr/JlRdvNlLceXodpr1yiapyq/
IQoS30V9bIsWxyt5Eg9hgUqJpPHS1WsaFLdsQ/DD4i35FJfBu08cySe6RldTHMixvBElUcFdFv+c
gdWbx2f1iU05l0TH2j0yRrgSc68UxT3rwl1ABKuRxdHooUTh4ypn8IR84RCg7Ix/yeJOeEg2Cuvp
CJdJxiNO/OiNBl5EiQKdwUrzXpahOV7R3i9O7vRWkcU3NXzM1RM2Xe3QJvyFP1qguxk0mbD1O+LC
5XXpcXIZWzbIMjjs45o8k/KUryw2Rbg6VtPmlL1yniy3qoA1Q01VqMdVMchCh7IEv1NHe059CcmQ
eH4+5uNSj+XvasfsT2KnDQpkP01nbAnVgscd/HTSR/GP1ZcVD/HmbypDBYJ56gBHP86m3yJzHhj5
7Ey2wLb1xPSD+hlQhZ8DWhRhT8lauWPL2zFimZTjYFcDFRzHyfFfdpTCdHwHKrn7a2M9vpu+nm+f
h5e5obwYHpKYX8MKYiL5aE/xK0fY1ql8BigIsgJTdzdJh5TERAQzzFq3VVKvcP9Es6h4zumy7129
bZ7jmlDNbZwU2KOtwMeK7oAbKbnLXE9DqxcpO/G3sexLRITax0nvbektUWzwFjZlXxv4hL1VURLw
VLVCSemtPtVXN23yYYDB0FgQu0ueRQ7aePLY5+WCTtCIbLWGlLCHXggs4nPujmXWIC/TWcAHn3c6
x1sFDXKNA54CUCnE5t7/XfK6vFA85ytY4WlBQ433SVuSgn0s7Ik0pVGJzE/48bc37yedN0W8GAK9
UYLggTWs6gd/xD+U+u6vF5a9rAtOwstabrPZZCm1DYX/H7QOu6kB13GtA3U85C6hkIsjE/81z9EM
7bRZiyv4k3UEvb52fRYmM/fbO/Sxiy4MooA2xeR3N3vFRe2Er0WfrhEuQtetDAtvOTic79Ahqtin
xgNcJEsCUdA5QU8s+drU0JleoDKEQCHcPV9M3UN3W284FUHy0XJmvTi8zedy10QVtK0ChbSRQuQ0
y+4fEU76nS174G8a24HxLs9ayOZWjlEM/KBLZwqtBOv5SQUmhbncg+JY+Jt4K726N8INrnoBSZl5
7AnvifZLW7MoLp2RmPo2eaE52x53kTVnvDOWO8Dw7NMJAIFSvUikh4xVSnmehXvkFoR6gk6L9p/C
ElDKJdTsqP1+zqTWHB6SNcO9D5khhzojV+8H/3BVtxW8WliqJT+TyDQ3BXKMxqr/j/vZYNSj1+aC
uOFKsR5Fo//M3MfKzPUGFLoCmO1OgoIU69vbIRRQ14jpU+/5oLYJ9SeclQhq9Uf20z8Nt9AHvR6L
NzM7hptl/dk0efBinrpykYkRG/ADWelWY9z5cXEosDL7gqgs1xWbO8qc7nWZ1YixNAZXwQQXiLFE
sVBS0kDvaFUoyjczZ0fReGjixqezudLTlZKlCe0ET6xLgkYpBSs/77abqNWuz6g4EHB/1RnjUOiY
Il4N8icdiLc1tgjYHFx9/oQ6kqWRyrkbNYlUKJ6XsMuxztiWXsYpvtPeAOc+K21l6/QHARCXEsJp
5U69HB14ou8wruomo/XWZLCFByEC9Th3TPN5eU77yR8fu0UxYRh/hsU7IbdwJU8uKpq/vnqM/VJp
Gu6geggDSFHD9KW22/wvryxDbmxMtpF0AYDamHu68FNU8Uahli+fXX1lXMpqshmDngYzIsacggdy
hI1jqhPYy7WdopR8msBJiFV4JX7QSRzRN3UEE/+BjjZNH7AysWAZL3e69zF5lYr2Lll8IRE7c58O
mTWAjndl0UkSBW5ii2ACaXUrAJ6bveINw5zaf+ntSAUj/SBpRaEdkZlyIW/60Y94adw/WrFsSLdP
tH9DQE6RrQ4B1A46wupCsgEFhTwmiqNaX8TACXxVe811/22Nk7ZIyw+CZrk4W9a3cm0yyRVFvD6P
goqjsRuOLBJs7Peo6hDF7S/iPnYrYKDssCL6otmKUyuUrwmWyQqYCuN7+pMhkP+dO/tjRfN3LP29
wT7hjONRx57RcGJcY5dO3d6pGs4AHySF+FdNkqL3JPqqFLpRRINxgP/6byO+DnDUtb63JtgJiy4S
ikOn5ohm3kQR86WqSlYuH05B61In9GrmEncCMlDL67vrVva63lZ5fgE6FZqpT2Pjpac6CerJiJuJ
q7F30req9XmeoAFwnlY/l7zs4rdo0JrvEk7sdPAO/mxB5Ec3Oq7ed/HGAr50kFydQijQjbWsVEgj
DGC9xfANpmzEnice7EgFQK2MxKs6UoZrbcINd85ZqYjjBFCD+nnikT/YPvEx6hkk1F8inxOhvWdR
20B1oOOzDxcjLY1ygauiBnlHDopB2t0DF+4fHFsYAOyueNevVdoJAVlnCRIZT9YrhybX8BM8RfRT
UVrVQ7PPNP7fvOtOf6mI2lIoFx77UGi7+/8PtiJKjbz2TUhwY8HDDTpiWeYQTn1VKTGLxo6XzZIZ
X5DSG0LxI5papzwWuCZiqhqijhaYY1Q9UUVVq2LE3yW34xvEDEf4OHvPo8gJWs7xpHVs1T6Rb0zF
igIoZ/oKjX1iMk1FsU5GIP+Ui0qqQ/PS/eq0uirN5pbgNboscZgQZHR/VeoSvmkTjhzQ4n3oTixP
pYqSmWCcz7SoOj2EcjbVxq6qTQObooTfZvYdDo4qMFomANB+ZGHb09Ol/vfVtSEnHgL4sy4AEce+
scc/4Iicd8+s+0P848BvNg0jrsf+ReSUcfvvz5FZZDJFtyWgDu3q8Gz9N2b7wz/9TKUhsYY/qiYX
JLi9Fnp46XSfEj6z6uBAekPl5GYGIireEMfv+CWMnH0++iYP5imgpzNUStaIerDVSPTrSxkE6pyx
x8ELY/wcJiry+VlASNc/iiDhDAatgH1mX/MANxy5WfGWpHQ/OMVg7CBCtIHV44ymF/Pmo9Gou+ux
soBEbDJrQvjrDTcanmwn+qFj/O8S89BVvtSU7AcWocK1PUkl5pGOKZR4wj3BONALRzpJArCLNwHH
dsKqeoWfBckVLXzJmn0XvOtzXWLEvB2ci96ZTe94jqMuaiYB1jpvy8INQkZxia6+NVuNAuPyyCCl
Z/6XHVI15qJMTqoLf3W2tohLXbdBXoOqqIX7fkiO1rocVjxuE4lCMVgxYcf2w0hkN8vQ6VNPPYpf
Mvjv/LKijUyohaOjcEI1NW4okcrpqPPIiOMPuJiiM9l9asoMiSFWeZLgq01IVX0Z0bVIPeE7Gcsd
mrlJ3Q1iWAAozrfUGMztaotDeFd8fRt5dWN99IOknRrJ3MxCr3tD/ZPxMKgpbq4pM2CsJxHKcb2i
T9tibcZ+A1QlJ5VZJnIXQY0D1ndW6FnI33W2K6S1+kkiNwRimBpbTsoRFVfDDu5FwYaV9ErkAtvw
Gp4gvVioZyPuRraaZmnO32Luv+Z478CxNKOxFPWHqc95ZYLQZls7/dKRjnY8Gd9lRssmYHESE36r
828a2tWRPe+QPGHQA22u1h+skzn+4Bh1Cpk9go7iA6WJDBO1Wd7RtGHwbb9ilr0RoaS1nTSMt43W
KXsSSVKC2aHGdC6f/0Todw8XNkD409VVamEafAGrl+/N9Xq91wCIAMEq7ARbV/NgdKx0KiFtjddM
juX6vbNu/y1KOWgZ27XRkXJ8pG+Q9v4rqEefpRANyljBsRkKaaL9NWTKTmQM6Mt6l4WwsBNy7xHe
VhObe/0vFPoDGXU7/isjE/h/yPKOY26JdyYnm8+6xfgO+ORwWKzbTBoUbapwyTk0x6+GZZYtP/fR
0r+jKGjAPq0PKDNl0B4z0bKoGyDKr2ZCXXTZVFj5DJmlZD6dkdCxNYAXKtRKNHy8VYMMQUJFY6Nw
8ZVFD2Vtif7jvw52WGo4A+++i1O9XLq3LMHieYSUnKYNf4zGle6m9QEu587RR+LRmKiIcFmpX/vW
3dfNApM+ORaCgbaRwBFa9jzXUMeggQKyLiibOMRRFaSGyUO6MJufacfz8FN9HRib9V5yQv5nK63K
SxmM0loIdDXnErZEJwUeCtG9xpUufIYNRRbA8ix/n0jO08kE9wKKtHOHrMgUNRmtTt2n1Y0fXcs0
H50dM04i1FhfXi/EiY48QCWhiQHd428Ht3C6nOdn6UVPE2UHnhpwjguOtjUaQv6bYc/9vMqQIS58
TJkaAcvwksstKjsGI1YFPyxOwF1bd/ur+JXI/yiKTrQakuZFcDlBQv+pPIX03scntw40bfG3PeQu
MKpd4xQtvFUOli+57ok02xt9omsBNbNhG/HurI6eqqT+pM5kmHL9wM2LpLzmQcRmbkZ9kQwYn06j
kDn6xu/0TVeNRlD4eJDqlwo4v4cbdW1+U73FvckmiiWCABufpsabK2DxKfKlOViFkPmG56qFLGva
Urz8G9gIl5uihozI+HimprAuNKEs3THN6We0nQG2rUb/ZaSSawcS/oiGg8xmDfUYV92jZzYJK9lj
U51PYbm9yEcz/xRP+gi2T2JyygVfDp4OP+aavoxSx2ry+5HzSbGXvuLtmpQ8YBtSx8uQAFciehBV
S65/+dCycLOnnxS7sJQ34cLmoNWdJqHBqjxrz6silB5nZcRMHaPUNQDw4a2gUQZmIoe+VycRbT4G
gIT8AO11S6y2e6hi3B+bVR4eyvYOdpQQUyPm6bIzo5U/hcEm9vnXc5dmliB0Z+PrN4nJS/qE666X
x+zEXk10h5nEJ3Wa5MRsezEq2pTHpvanK4C3FvXt7Wt01x9pMgaO3W3g8svHAfJAeSzPPrmsLoJv
PZdnmDnOniggu11EOGgFiWeuoZ1/2U6hm/sXPQfr+HV2KHwsoxkO6+/TQMC9eMqRJVNumuWQA5nn
O2cTw/VRvCLPYuDoiHUy5RCF4/mFtyTHqdEg3jD4fSzcpcpBHpPl3KBhEa+SMw3YVRctmWdu9PI5
B7fGh9Qanx6XtBFqW9ZWwJlpiHSYl2ubVxr8F26OfKVS3IOEAjH7IFQN+ihJ8dkpQf5xFpS/3ATL
wvakQaXQJJ663LjnGd5P9rzPQ+l0oKXHj5Aa++fWP0xnUQwpr4YZN9DPcS9BTs0lHpjgJ7En8OYS
tFv6HcgOSD5DCLzvZQey0aCOZ+aj9oaN/ZXqc6zsl5rjMltVHXtmCdWvtPQq6HI129+0NjdZj8Je
7sjzViR1F7d7MTM0bjBsokIVr5GbRjtBGUTf3MuGu9Gzn+DjO9Cz0SXxb7Sr3h/LCa3Emx5/lAcD
6SR+HAjt+IEZwZ5L6dPDh11hDsaiy7LJBI+EEwXJ5tTDui2R3iXK+js7ITSRk3mfSjjcC46IEuWs
e+0zRMiv1LVoKgh5ckH3b5DZTbb2TUASiLWci0YYT0vPz8AJQYML4KJeNKhcK8ohOvmdyUx+TUjD
GCmkB7i0n7TFNLJDtaLPIMjt6Ak9XbIvU1Gql3nHhFuvJ5q6iA6ToUN7xG8bCFJuJZwDPq3lV2IB
xs6/xTMBKziAsJ4YSFBC+m0oc26hxRxKCdwF/YBdIBDAoNkqYpIdD8TLZixSncDkos5GOrlxZi2j
VaFUfTp++hZpipinsjJlDqX8TQakRyQSsVmTm/VgdaJkFe3TF/lkw1P3V/6e2BLm6lI/6OQPQtuS
eGiXhETBJn33sCLRyO1rDU09MKqAg0tYoNCutXI2g1O0Aa7QtgIKGjEX/myRxBtJHoMDKBpNuSLs
jx2CfeKXz61aQGe1a2Gb9S/xAzPJ18LBXUoaSuzFPv84EWyClGAAx2foJJc9ZDaw5f6wbsWE8O2T
7JHh25XF5Vsxem57xmVkipM+nhjXyRzL8Agpr/m8UMETM6UyCaCLWloDJFwlcbyt85FLLmYGUKvJ
V0cfPmleUTc2JRtTr6G0fcy3GGs7+/bPQhqvAxJYJ/ABENCDRj7Q/T81So+lVQG7OuHhI0dMcrtb
1i2+JtqjSN3IBHkJTUEcW+XqF4wrKkhEVjzpiDUs8m95uXWdooM1yd5UzQNYNnen53yekL6OOMdh
bHIiz0BDDF1o4K7PcnsMpmPjgDyVt065dnNvRuV8xhssNZfR6fn3AWqG91P4xkD2C+jmcmvP4hXP
AafcBgWlizXqb1mtKSmKNCzFrFxsPBeSbLCz6p4s+QoplQxF/82eZm924Zrh639Bl2YiVPq7VNbj
3Amha7hnD2l7Cl9rpuvVrN4XqiFIhyGu69H/ebbBz77uq2a08kQk/rqgb+Pa4sHhyaQ+IjNRaM6p
ieeVAt1tKPHMRQUma19evFc7odyFK61nXEyFB0nps8ZHUCWQ9Cof+J4cMtD633yb+M9UdOOdgeQk
BYz14wGYljp4vQuE+nrrS1Ck1oa96ZURu6SsOjK7Tko2EORoFvShtZdyscG+1GgYCLeFJkHvXP75
O80q1MaNXVCUB22ss/zp4Jo2PDUVH7vfL+ztbyGm/4dKqKvwgDerz+ZjqT5fb8VW94ulQdxwcucB
tNbe6gka/735iMRAdCnpIatXGf0A2FgyBnBIUD2CfYmJti6ZyIieWmf6wnYFg6J6iPY8BeUOJ3uz
JAXLDiZzfKVwFjyxc/v2e7IvZ+6rJU2bYDqW5q24rNpVkr3nZWxS+sjvUw+DisZjm/e4Y84mkHi6
PA2pykYhXVKSIcpZKNgY/ltHaM15R00v6qq6VFPPzB1YKhN5T+lFPDRt6LtCsKGMEbiX3iuWGb0y
gnimGwUcSk7CQ9cA/ywj38l9WNIhzB78e9pHiMJmZfNaofOGXfpVxJWr4UAo7M953lX3zho+5qt0
jEgHQAKGWZ+ZXrOPM77GUDVEUydJec4lOypdx2kaTdKAmQ5pVDbWQV3iQQG98K6LNMwX4Y6/7Zf1
Nd/tghz/i15rcPQUL8JbKc1/otoL2CtYfjvAwhEO1Vzo19QOFb7gI2szKCqMCNcu8dx8nnStMRuQ
D0iWi2mPGbyLDfZaXMrW7SwRUmup86BIX2YtMDO/t31t/GgydInG1kmKw3Rp+YYF3Iq4BdnJFE2p
Wjw8imqGbL7oQN4NiPBbTcU4VQz8CG7aNxkAPUv5PmF+G4K7QMlwERaGQxrqbxuVZ37rkORU/v9C
hPIKDZj9pu5/wuLHp9Ssv3/RSKY49cvm8CW+r4FKBlzCr8m/6FSDJbKrMtajx5cGxZZ207ONCfnm
6bo1dwpvTl3oLDcj+7aVi+DOa2XH9sDnzjjNMhNpitHwQEEqiXdDvsqJp5Rd6Xks6j/b+8KWudLs
Y2lpHPm808CpK6rx6WATli13A7yDdQbrAG8qeRfdaZDh4aZHBxYuM0pQUzHJfHnxx0ex0oawCXe1
wNCUbMOcha9el2046ZEGQXGR307tgM/2slVJMt+kyB1eiqdtgOUcuPi5Gy1jXOa3xb2Et+mfW97f
4RFz98J8QdV9y5XEmPoZW8tSn6VS7lV7r3MZrksCmYx3pM7WWohXGogm3GTjQPKwZOW744GcQOCz
82HZB2wghed5/IZjJP3t3mdeYwzvZUGeS55niFuHgjOjwJhLABOHO1jd7e5BQZn7OXIiNjxNYGZy
W97nQurD1zk1LkftL7w6YZqYHt2V8jeZS2e3fRXshAbZWdjXjIbanQmZoUMhIGUlNZ3DJxvRIYxj
3hYB7xEKWoz4Hug7zvcOVjCluIKWSA4HZSlI0VCdVXRa1qMt5WpURWZtyYnCbkpPfOWRtEmR8V0P
nPXdSq+YjzDlEgXlOkWK/hfYw3v2fflhvh3TblpjveMGIkeFY7mwvJQe7359RUeMbImRrndYm40h
g1NtHmClDZo+psrLB4dtX0Fc56veslfqiel7jppuak6lvENSa0xmrOt+MZ0X2KCqQf6s8Gr5I4hR
fNfymvCycHsDxU6EuTZUpmCUgCzIdo9ekxXVL3Zje5bDIDiVB+f18x0oHJENwU24W1zI+HbhFBjG
+kC42owu9RBEOz+jw8gvb9Q58/konCvl2PjOYrTTRqS9U0AOHs7BlxThHN1HClTL3WToPiMhOQGp
xX9iermXxqI/sK72gHnZJToABcuYZDRxJJchNtQBs8dHwb81iG8apip2PyRYaGNyIWIa/bFj4Z74
p34AsSfle9Txk1LbYt8J86sN/9zxpK9if2jqztYtVRs6QVjMKZiiRw+MstKfziMGeba0sk92Ub+4
y904Kcn2W5cAsvX0GdF6GqJPCHXUyq76eyCl4P7fnVSAemlQi9VMu6MgsGshH2/SH83aD6P+bIif
2IVgalpySInBh+L8+5WOVbwXi0+HyGfWpSWqToeBMPT+eVb2Kp/pklF3J7wMS3CEHuITvC466ehX
1m+vsLRTDEVI3w8hksVKjIwdMDrCgrDa+tmyhihMnEU6I/oeIhHY8YLsWQdK1oJrsYVVmcQKxdYI
oD0jAJxZfiYm+bo+H4h/0SvKawVld0UN5gaIQEWTPX/ZYBhciF7vKPQ359lm9ZtHK3FjN/Lq08YA
lT/pcOe4gSPKA3B7BJVxrgukaTId4CtpS0NpX2L4IabOeipgrc8bz11rdAOkcucMJzScJMpkBJAt
I4t3yvGJM8nZs3/iGrtjUxHSEZcb/Hsm15bmDdgmFCM49XAs33XfVAC7yaOz/xyzcjXLCgpkA6VW
LjfPQTAkbf1vp5/IFGjNGB6axhLbU4ZCED9BQC2Rct6us7iJD4CTadqw/gZ3IPS/d4wJVrEI1buz
ssjprIBGksvAf7p6q2XzPV4srDf3/h9egwK4cS27346mVUzgjOOlMmW/x3ejmhDtxUDVOl9AnvaQ
K2p/Q9d0YfuRFnXd5olNrJkSUh0C76sya8Ius/zDOVvr/oaJnf61N0r+smtpGjZMXBYOxKOv8RA+
3TOaF9szw676zlat1yPrDqtzvS9UaPBhBwouGH4Ibp9E8MQbcDvvebZKVmomZmlOJWN1CqYJ0WCh
FXem0pPa/aioLvco5c2vpSU7ulD5ekoZVykqVpN1zW33qohjJWih8Cxef4salOLGjFPnTAH/mQBb
BVA0d42m06vKDRCRllo3XpAXzRBG0hXcJZ1oVwJZKuOdyGjmiQtYBsj4ceoMw9EygAeURC2vvjgu
9FsYX1slyD2TbkmrcTPlkI5P4t6s8RBRRHwh2fLSCYEQoZ16bDj8n1mgKUe/RULYtdlx8y7YKfRJ
V6MnNgO5JpkumFnEkmQy26iYXGuroU3CcrHJKr+eV/3ugXgg/vyRlHewGF2oRW1t84YkcQqdiq1+
TCMw2J77rA7lYcI9ke6JWmp2bOegyLc/bSerwgkCM2GCVDJ4E+xUMFwXPuGXoyxXSqIv+/KYl7FD
gLjAlorvPuTqJ9pKz53743CFoJYPyRMew7J+iFI7nvP6aUugrgO/7eWmavoxBYuYEhMqcBl26Q3V
sK6MhZRRBrTBPmDucUBUI75YR1fFMlsfifwg3T/SkMqv5dIVa5g2avKg/Z6FVwM2UT2bKXILw/Ao
qo9f0qPrcybDRluOIn2IHclfSDggEXuGbxle/a15INdgHGoC2wpu9rXT99lZNcq3VBNOwlUsS8zO
u40a0ka54S2Uk1XeA1I57GiaykgT89c0qJ8QTI13GOvUkMRQ5dVTQgD2EKlc6X8wyxtNd1lZCGR2
/XSNLPTrH1PiU1c3nTpX1DkfiXXeNRCGkrASgHGYM/kjQULeOM1SLGuf+hBFLm9vY3a/w73njBjU
cRZjDNQ+Ou1kcqWMEOgDVMjg7H3aFMIb0nESO9VrPaEwhASmGah59bbknBn0G6cqZmQqOVBhdGVt
1C+HdZvnGQ332yL9uGnoXA18vavIWUJVLrCWW7iQ3/7oceTb6zmOx6rmH0oCKj5zYXg6SUD0gTfG
V8KqaYv9njHkWEvkzxuVQ8k+mqJMhLigTM2ginkyzSxKZz6FmdLvlq+A/P8gVohGQPw7Pb3xnJn/
9z+XygyTk6B3f6YSqykc2WN1H5y/fzB/QLTIpLQaN1sDsDeyi4UoRAfknABoq5wcZ9+NOd4cn5L4
hv9ZFr31LIfgvb270BCZh7xbEH3gd5hhqBC86nlhC6UIUsvxNd8bsu/nxWHxR2BZLhsWvbNHB6IB
RM4/hbf4K7m4G6wmaFuSWoOLs4MmG5MqdBJ01knWMKpY3E+rgfYYN/pHa1VCJtrD50cuXM1OSkLl
jwuRZYPfE+7Mo8HyobIbySJV3feLSJOHWGgmI3jK0C1v5k8AJNOBU/HgRPEOMGfKFcs6aZkeYNwH
O7+rzSXRGt2Fu8VpJ3hQ/w3op2z2VbSmSkND/zx9MxcR9wEDkIagtqX8p5GAYQicp/IxYLS1QQu1
i6SGv2VjND6w1rEFZ4w1c5vZ+4RKyG/IY2Vks/qvqfcAiKJUlhM3rr7hvjV2sJWZkmJqPzRxHdnb
1c9fkG53jPtoCeaJpe8Rw8FUYwxllHwYnVKBMMO0P+f/eYnUYFBsLQFhsZVJl3x6hvJzxshBBCgd
GY/ODXrYnlLmsq5o3Gkcd3kNx2lE0P17MDhvZOiWSdpWYZ0/1/nNJliA+38s2Oh99BcgTQ2soFOa
mePfneAi9eW2KZirdoqPjSeqkJbJ2c/HHkZKrR+qxMG6uZQIEzxRCoAZwAgk5/5C/rQYZt8rOYa9
b9LemI6CZi+MPe1+TMHftqIkVvuOOyRnKMtJpggw7m+bM/cGqTkqPKwPHr6pf0b49T4TJD4cjt88
SiM2ZQhQoV9b30IavdWcplEfahOVcDvrVFju5dOvZp9lTUdw57zeEE+yaOnCH+YalZrvEyulcNpT
AyeRSTr3S5dwFMupeV5WCQQJJDtKCE9C/YklrlQZvxGydpspt3gRG/xI7wgq4nlJi6lFO0SiCS7y
SSE8QWQavyGn016Pd4eZVJj0o5H05SNNWchXPTdo6N1I43PjwYFLEg4kYPtBkksbkwpj7IBxm8ov
03pMJ+OZRwe+B1Q1MPFPOs9o9LiwXpGRNP4bqdsakD2vfKKp8yTkzzKwceSfqwFOHniexTEt9Ulo
OG8TJqaeW+7tmo+Yyd1H7eftKfsRmTygSnwnRDgNnoll9/HGx3jj08qursPlARP76BYorv9NgD6N
SM/ISeCGR4o7B2vKLG2MlnBJVLIIE4rATz7WQLCVujGsqG0V9IHAVgEfg+/WPDeKx6nVVyNY8AgI
rFM0LAqniOC+H4Fj4ASE3FiSQQQNH7EUXInJfDho0GZj7nlik6oL6snptydj0BzQVzQZzj4H7kIL
JWEM6cvOXrOyJA86HJcLEUFF04MKV9Cyudopitby0YC7kT3uWwPSK/uc6b9VwwM0OzWWrUXAXeRh
+YZJFNtx3t3RMotV/mWuKdjRp82Yk9ZRMipc4cy8xBzK2K1PqbuGFjwiEy7F2ipi4gavyXq/cO6X
S9ycSPkDbR28J2OhBu5iTLyM3xfZ547JLwuK68PNDnHU5fb1/csS7Mwj9bqtOLZABg8XtCvGQBv0
cOUNXUBeNj7/rBfgIMei4Locmlls+iF1xKE2uIt83S/xbErxQNW9YkDQjJa/CW0kKd0YwnSW98AJ
0/ONzgfRqT3DElVKha88SRUo+AQ3PecA2Ge1OL6M06RC34LxYeJwM+bPxbI/CBzg/ClB7CSSkCbU
oDf+KjJAyG6BzCBqDZt/TMlJakWNPj68OVMcvPVWUnt4EJ/FTxkVKK3VUFYiv5Xrnm3QfNxxW0hd
xZxI74SfoxxMeubC4ssX4rGIPUcuNfsLbQDg5T0di82e5kL94SlWTxQg0naYUiQGq/D1Tck/dMnp
xJYqnnSzPfUyR1TdIbP8CreIj423FaHNGfZejIpphxXaPOmk0PUo5eN9eXINOSL23BwKbfULRDZj
69I6DLlxV1fYBNPP18pRv6OVOKXoUt3mwZzzvKiWqe86QzO5U70gl45Oh5aEm04aGzmZxWB1D2Ez
XNaYIwNlVhHB9I/8xpNU0fY2VuMZKmaf4cbCSd4lBcbCtORElTVU10M+7zdn0MK+COjPK3Qeb8X8
O+hthiV6REV24uFBfLhUmEULhn04+Z4q9+ldj6jx2Q/41081yGDYLHhTrWzsOX5MGBQN+r5RHOEC
RiD/yAmz57lnLmQkKmEYwmJZAKRGtgKVtiyOQX6qA6VWp1hRIfMXWJYeySqWLMwwxLR8NEhlKKdu
TwL3Cx9iwZ7brm2mRUAC3BbAr1doa74SEnmVEuL92H1/1tHV/kmpAeRHTazq4oa0ASI0loLkJuJS
fwbRKdcFI5eBDXDSEXDjvnnZNppqdVTsIDR9rZiSj1CIGJTRNHQDVy7wjqhAvk2euTctC0Qm5EQD
gGzEZD5P9P1aYy6CiWW0ZV/mvH++zX7iRxOaqZs6Rrud5dH7KAFdVy23FiPgzahqJ/y4m1u0mCtV
kTWCHCUwcrBrsFY8J8U+mxQgIGlV3vbexon+7Jz7CIz6UUSXh0b7I4Dac8NX9KvnZVC3X4hPEgoB
fBIW6jNfpL9m/MmcWwPYUVcXHYsedz3Qk1YVVOjmGs+qcXMAgTONSxtzGLQ1+H6A6HxC+gWDdXBo
xURW0qcOuo7UFqerxPPjROLo3OvjUHCeqjkbcMuc/sISc8yLb/NmoFvYtrfn/EKMLBIyrVl8GEtB
E1+63+a5BR67aiz0ByAWT0G3qCNmRot/1gFDG9DM54/qr2MePN1ubUsYWoI+FcXaFb4vaW326fzD
NbQBzyrmitFcUhckxmQUvagiTkMeekHiL6RaumrtbGte1mdcJwCSq2u6qxeCinhY6CuiRPQ5SYIl
RmsLy7Nb9Fm6LdX0wMeGjqDCJWYBGwZlhtjwU9aZ9HM20Z9TGAilOSmJ5dnp3fGIOV2p2O99pnLM
f6tc6Qt0uJYJQeYk7o728ufPRt4ErS/3tUJWwsieN7KZzjUO9M6Havz2nqdNKNrngTF1C/SQka5V
JDKnl1ygfpk1lrQRpBmVrhtdtp+QE/AV4/LqRhaaAkRy36ZCwyAxkfBaKY+iC05gSKAnxECTtaoo
h31DFmB+XcTK9ZEKjS6thkwnQwTERtH3UkOKSQUkQ5uguMf33zKqtuTawXJXiu1uNJ9ZBjNMM6yP
E/vueIermF1MtlclXHSjFeg7ik8Jj+fiK2qbAogEcwglpNmRwFlRZ4pm7MYbcNJXPifrIH4BF5YS
1f++g1HS5JkNuDDECfFNApEPYGhqNymErOQ8Mp0UVEcXehUA2vItmvo7Uo90fJLD8KACUiVjJkNa
oAlRqlNyYwHQVBfQITX2zfROOa2RZ5HqluJ+bXHJmdJ/iXzUdtFo+bg0jPItNGyWEAniRshEIQq7
XZ8h3oD9VtiNTlCosHxii4dtwipYlGCF+7C21hnu2YMj55f89fHHdIMydtfNMkyVhmpUjrk2H08O
LdUNHxD/3JD6DX2LFfcDS6RMppfz7JfLr8jMfprJ3VARU0WeD0zeqOxKctaNOLWChD5aJFkOfL1z
DhSBZcRjFAT+6U1ZyW8CpC9twEKPv9RogGA26Zzm9fSGAre9F8698NJzYSZln0Okk/pYgaePBwN2
x2eXprxdeZtDiKjD3LtUPCFDCXvpW/UNg0ru1bGy7higjzRrCx9qJwXjZg16xYEeSSHQIWb/VTjU
suFWiTP6V6pMD006S/IooyIIOkiknrI0ndnSwfmeJkMX4EIgqJ9bTHRSY54bHEErooQa8uBXmVh/
9/7ZR3t/bwkhgMJdp+wKG9AfAc22Kc+ILQqWbxxF9Gu5a0mQSSjf4E/YgSNlC64yzs7eXgrHHN+X
XHAMY3q0Tk9xk20ZoichbGII9brCnUmjjj2MzyULSPtafOWoFS0sGza5GoS0gS67ZT5spT9zGbzj
aFabZztdATsTk+YXjyKHDr7Gs9u8AbAYFeSQcVCbzztdqCMX8whHKaMWLMK5/h+RTWDGVttdrjno
N+TW+nIaRRz9TzJT+lhw2XdFWbYATPMbhPcmudbgiUvcwaZsv1cvl1ecGppSngXL5QclUzRSnXX8
O1nJPl9jc591vI3/orr2+EVVY8RFikxpFAU+z/ROF9H9Kgh+I5AOrQZF4P7tiaQfIX9pjEMcMtMW
wQ0G6golHvZhqVLnVht8C6z7tCNzHQ6mKG9/XexHbkETkx/j+OjawXdqJfn5U+73Uf1SE7a6KmkZ
UfmCadZiE2zmRMQHPh9dT9jc8oB1NFdn7XTFROOhjWuELhxvDLo2nPh84b72K92bzZ4XShFjBMBE
Hg8JeE1RZXHd1AKuXgJDDOdfLaku5Mk/ACcNAMNwzHldvkEmDkArksNZfdEMi3oQOyacCTxqDo4S
t9zojLhOiNqG4OY6k56oqipjSGHUYJqyrMYZnkAwcYMp6vzaLlfLO2Ty6ejf8r/0blp03H6prx1L
6YUxrbPG0ygR/MwHWlAzYoj5a1aBqenbZw4aZM+xBkmc/XQEq3EanLAhInRz9BwogM7+jggr8U2g
+d6kVp8ZQxx9tQvJ+TwmeRaEeaqZlTTIfWti+XPxBLq0NLdhEyODvg1E22wXL3uzfOW+2QkHSiI8
H5SmeJlmuJbQMolb8aiFWBEUdY+ZNg/LKTG2RGb17eumFhON7oVzLs6TvdkyCQBg6tn/I+BedMBD
jCzs+P6YBBB4OdnGZCHwUh9Or3QYWU0hXDNfpT5v6quyum+Bq9hDDxhDp1RSEhoq2xFZ18+R5Qjp
nxUs9D3fx5woJGmE0MHstD9YMR7xDUBnlCVWEoSW88loNVTXJGh34J72PodlM0tMsLUN0MeRE9Vv
i4Lv2pU0xMr7nPKv4kx4psjQhG5MiK9o9Fi66v2rcxNGpwaJGTUZB0h46agIY4LkMFXhRpZJ0kHO
X1pBPG+iK4CnrDQ4EBSV4JsqbD9T5bt87C4PVGZXJIUmrq7LIiMvGCWBuPWPoDwo/UEVSbmkR6SE
65+3ZHIhLARxkkBAnWcR3Hrl1jQY1lPqZz3w61Y2u5f5/N+J/afSxr+AFUlEIkTg7RzOgU5Ul/tq
WUXsHtzXc+eY5jsrYW64LYLLbOrYmVXVKj97wulOJATOs0KrTo1/RxPzJ5VY2GQIqp4zDglPu0Oh
GUy6ZpeOux34GiFis3jIV442qLkZ6By5QaIZl+Fvts+RmIfavGxpe8UIOftQqkCZ7xuU2+ehUPvb
r4unbbpJSYScPBzVhhO4qX4IcZx199VCOKDMFCOrn2KJmdZXQuN0TyoM+7mRO7KUVGxdgQw5cspU
5AFXcSa7AfKjlL929jiXtGojG/EKxb7i8lgLg1xpw6I8qdukRj6CGT5HdSnkMD22nLOLpXzAn4nP
9UwGWWDEl4bKY7Axs9ZOna5BwIMFb0b/2u3EPhkjpEkmxf5p44P5I2MidWYIt+j3I7bdbRIk0Z6x
/xjrRON/8Gg2j7gkYCQ1ul/oBvLRPmShUkRs77ykVf0rRvCYcpu37QXVGqtjxiOaCXWVM2xeP0/t
ymYHBQr4jOeAzu2GhV7uoJfG9gTNKh+cobW8/IxONi4tGVgF1WaCO80enbisa+PYBiwxqfYZcqYt
XC22uQe9AWSi17EmhmaCw1af0eqzksCJBlF+XzzISbq1gf8zT88YLdDg6KC3XTTHMbN5oIfTDsu6
1P0nvHlvs+t9iX6kwQ0Y6nbX43s5K8B7FDwu33fhzJdvnzCBWpbs5JXsBNs4I/EFffxm2X4VxchY
1J80yluMm5ZwG98bhO1qKWOtN1GMQXQrQDTcvQHXcTuR5Z8viU2ykYwFY1bny/6ITqiYWcgPbvBj
9N6cTHcoJ8QAGq8RP6/CpM8JuPcRFAjTmWOtokYa17ANCcBueGaJTH9wpYJcn9sZtWJA1Ya+LVnQ
5WYMllMgz3CPCeXVueXqEUWYXYCuKvkZ1dvyq584ttOAttIb7t82vxI0ycKLuf7RZjz8aTw3Tfkp
bQol6pth83Q0ug5OantgtO0/37zYlnViypA46tb7Jp8lnHr4KqwfKoMQ7e1cCYQbDHJy83BGRg/O
U2d4cFaCPJtz5mFZnzfbkXiYDKRmvjNbctVtrARJG3OPtZnDSuxJMnNwVlV7JEu3PL0No4XhH1Qz
DtLB596xUp2KwZ4R7Rkc+PYWXQ87Wd9jQpfsT6u0MzkBKYOS9/ZedD9kpZGtASGEI3F9To+CGwRT
AiB/CD9sWE85XcbTVPUaysdATGmEG8E0VUh1TBdwAwf92JlBsECCbG07DmOxMpe4e4vekilAvlWM
5ImgpzPqJgYbbANzS9X6ZchANRfNcgQQ2cBUOJxu0Qm+YBTlC11yuBiCKihMvaoILiTzTuf1Nr32
uymPnUnK/i4WZHkZ7bJZ7gfVWhcNr2W6K0gqmLL43+oZjX46lPnHLOzafOLgW3PCJc6niVCyzz2B
ABYbwUUkt4tgtXum0AuzZ1epeLGa/RksUfkKt1SHwtuEOGbJkUmkBliF40KFxc/Xzz65stwZgP19
m8oX873z33b4MaTJqDC/BhvRuBCGXmVbyS18IKt511zKMuUX99RYkrWIiwgXwQRJ3wTlXflTn4Zh
2xdrfglnvajnNNAI0A3KPkbAzCbbzXl11qMFsBU+X0Lfv+Gffr30nWGIwGm2bCE5E1peiOXlTs3j
Qg0YDopPcEMztb/BNdhF8DxbV13ksXBdQLFe4oqSTFbjxejU3GEDHfAEDZuhf7e/fugnWir3EvYa
35M2pDhxxXZzNFTPGLLtG8LOZ7QiFndoSltB8f+dwC/M9Nodsv5PgPdGeQvnapty5RbKsZraO4TS
FWrZE+BptcLISMipswgNMsE5sNqZs+7QecQm3+h15ooWjTp2WTCo7S2eY7S/YgedXKMvw8vEM1AW
UOOMDLBTQN/AZA5p4WtxvkDZcL53oh6jtjSLkAzmuKgwBmx9nHl+LhvNiUcWbeEEkEqZ38xztuyi
ggfCPADUQaD3XKe/CBUKQLj/D9aRyofgjJr3GX/iuuWZ1TRHaeQU79cRrz6Wdfcdp0E231ypP2Bu
YEQceW/j4NoO1RI0vYRoeri4Zsh+i9HqSQrCJNHdUrM/7zs4TG7VJpgZe+Ew+IuWhfVRTVh8jPOt
AXfcxsqCv4GbiPLjdu8pFRnxVwEeGJFgawLs5WqrhnzSS17PfXpsJVYeUKJajzF1eU9nSv+oH3RT
R7SEW51gvpQnBcxBuREDAytJlEUlVtu/8cTGr1MQhpdYH9wJGCYFkHkwuWFtbvXpZr9JzMZpJeJL
k3FWMTmacvdrfi/ky+rB7tfwuk9IhAVZg5PZy+mI/+lKokr/tu3P/Y06Znv4wZmCRoaUAq/So6HN
ykW2TuuyS9fIzJY0sRccI0vCQTerGror0BctACryNK8yjfai18zJEHTGeU8NCaQ2n9KacLQwhFRV
abwkNqPIdx3JBZXzUuRFUEfyB2b6wE584AKpD7pF16ml7/opW3t7iOjM60U5tDXDxcyn2f5oseaV
Nj5iyfsBRyHCTTbXOcN0/PKeu9tJeSiOiQvdtoxIYIAC4tphiSZ7DApBnmc2ZXd96SNVMkijgaFe
rekWhUMkYPxZSok67r53qPTxgNo5OjaQUESgkRadWZKi0zI/Pch5eWEAN/kE1FCVv8P4pQPL/Rcs
ueb0A6OzyTUYL8PClnYKMqyHJPgHzN05hzEzNAt/IJWzbK/CNu1/X3nIYMwBRguVPd9B9t1wmDZa
Kh3U96aBtSpP7br0y29Qbxa9cc5qgkqTAah6teVpiTCZrWL1H3vxCuPxF7xw6NnAnWEjB5grWyV6
j20Dv5v7cz2T7R3omxbcWhHDUzj7hq065C3QXmKwbVGuiRDfDARn3UXgiUBJ8yBAuL4WlozhOTRz
Tzph0H7zsWF0HfCJB2hU/CGNrL+HBR1foB/ey9qOoMIpuGg8BSPWiR/E8Ws8WzprxNm6BuVUTWeE
QKI5w3stfhDs5YXpQi8w3OXP/z8SVpLMk7CZ4jxnWFaPjtJusTKzZHrFIhpvEb3pN8QnfC4ilj1z
c2Dz1mFOvmqryJ0bLNWrAnFP2NRoluBumv4UtxGPrrulf5VWpEJfXoXT3U9RxR8x4kwHYjdD+Z4D
x5Mc8XfKorxZB2a0iX8buFFTohf5Z8A8KgdnZRzvDm9mDLlSSbX1zJtcZRkomDnjxrascf/sli++
3pPEDpuBaOPStIxqXsRuGkSZ+oJYZXRDOtrJSTid+/d97crIAE6j0kZFUU4PkKt3i/nD4EG3vNWq
AvnZxmMcCaqLvS7qZZqYa6WQ/y/Dx2jgprXC/C8ixfkXOYnc3+lQIlIzj6JbfxTAsS+RzpYjy27X
ktsvSBKmwkheA+duSro6PVT2uiU59YXWP+cHZ5S+/oKKJwkll2X5c4dSqCE8p0MN6X+Y5nXne/Sg
CNoDO0PIJUwsdyY5LZC4nR12oDDcKV81MMyV3MhrvXXOIxS9oTDrrnIzE/iEaEXaqAMenPVWxwLb
ei9UMIzIrCYeMx8nKbReF0VwKcgFRANpfy0Y00bTowkiG/ygIRFy3mgfY6YJvi3tgcRO4RzmffsI
N/eIh3eD2sqyV/KRRu10jAJQfS05l9jcbeMECUg/vH8UuMbbMCCjpxSuWo5bmW1Ve8xM6gBoK+ht
PDFIqRIBXGgNt91Xq76sv+4DO6S1UKfrWd/nH0a5WU+NScXB4JDZirCj+X2Wmeh58XS1XZ2VhRhW
+Z1aBOXl+KmZlGVN9KAoHb/2B0z1zTKKZyEf2iX/+P7wSSbRIbN9AS4LsYcd+Zzeoxsmj4ypZCnR
a6fB5sU+Hf0n25qtTTveU5VQuT+Xj1JgyA/MYrMna1BUDdCqUy+yMV4BF0SZ26cVtnSnz6ShBoaD
nHhpgCZd6ZjUxoTWmMZPjAPU++O/fG29LmUu7LqIisEf+lNL9XjcDqE9uFP6eFKZ4x9jePtR5dua
x/EYJFTx9rPNmHs+HMZI30BNYp5ZeV/XTgfBC0kzqL0Q/CH1MBTKi7vE3GMyD3e20x1lYgm9wREO
Zyxp5JaAHdufsMZ24WGIrf3xw3h5TwUBZWi840jhNZInJ+ha85VmdSbLtGpdJ/YKochUeJY3N+AW
KslYVtrIfHHU6zauoFV8nXvCOavti7ObVYvq99iZ2z2PZnebiglzrknqKCr0W7doB6sZ3ZajUmb1
TpHd4EyEHUIOQfoptdnuDGWml/uxJ2OJzs5NJTK2IEi8f7rYmpjEolP9oomFRpU4WoOHwL96Nk7f
WuLS6mNtjbu5kAiYMUttfROdrKdCVRTAm0NVkIendAM+axi3XPb1g6+3T+sD2/nRXq0B6KWnrPtO
4ZjkN2sP38gL9Eqiy3jKr1F12+ozn26S5psRUg2k6nsTHLrLiuSVTwBlW0ZkR7XwpU9NCGtfwtY4
2QVpDCexmWUsV2wDa27s5NVqo632nY7kNxcrn4319r6gCvGYDQMfYhYpB38qOZnJCgzGrpbgA7R9
lbChKTElCulEb9ajv2za0OxvvJdRaAzBc8iwpvmfqDrWzrHsBwRVil/44fHpC5Q5bBTFRi2STOXL
5wqHFzpFwibyoWr+hD+GB9Q0o3675Lvz0w87ccWvylGe9+KGfBPm59I1u1kiWNFZxNs0/s5BgM8B
MjXNTuDYuF824XAUjnZCs7lbm+9jw1HckH+SXnbDJHTYbnrMbLpF1hEHO9qwLZfZesRhvwlZFx9n
KiSzdvnA/VyJOn5Eo3+Zkg9PEj27Ylbn7Z6HyfqFqN5V7R54PeIRrHhEbxQDCIwEtfcKjEkU15NI
fj1cBvZYsYIjQ3bZD81+gdLxb7s9JYKsdSWvzFMH7znWrmrp2VX7BA7LaHLpohxAhvYge/FBAK7u
lGE9+0IrIuvAjiil5vWGGqnaHLQY9+U8mk1xkzjGw0CtiCvKBXNpl65PPgCkVSKZfPunHlXuxGGR
jGqGU+wKUzHmETynHC068eI+AGGn7mzK5TQ/aCmJ30CjYu+nNLpd82qk/Zy8YQ/GXcDBTl/VCZhr
WNavlXkvKrE0sBKzO2uIcSnB3Vko7CD43LLUkkj3Bc2LM614wXoNUqZXLb18F/8ZmYF0ogSHAzc6
rwunX5YYKavJffkyhOGJ8eutQ/w969VJeMaG2801WbA2guLcyS8GxXJmCFX6F73k8Aw35cJYR0jN
cb2k+N8gPZ1ca7qrtlCvDD8mcpa7t34lpHU51Hr9fY8yr0ZHKXRTpKApGtF/i9NAEUa/Z3WCgphB
aa/Vx9ooN9GzKXelg0LzcHFFcFIGnY4dF/PUCAVOPI6VbSpd/Nk0I3DTk+0LZVwhZa4BSMVAKdpK
FuijGICTsmT8l0HuzWLgGLjIPXTGCdvAFIvj5FQEVQu2Viha4CBHcVcQS6gMrban3SN3dcW984K5
nrG/vVLzOpqYFGE5yfIpM6hHQI5m6YTZZZHUi53/NyWo1Ped5BTje12xEO7wmy8DPZIlMdJC/0fk
sRkSUCpU6Qvz2ZLeLpbFv+gLMcBDOsdDAbU/eHPe8heEuJ0hU/V+T0kK3Pjb+QSBJ/EW+SX5FoUd
Wsbrb6kp4vuH3/wZm1nH/Y+owZVfHhvAmusRiWhVo53zC64jXjI1yAwYHoxmuDl8Qntw9GLdb/X0
ICTCAXqqiv2EmDBi9SnV7Itcskx1wC8GP7OrxNqNi1p8eVDcxY4+P35SmTt4RN59sJVB5sKN8i2T
uP2d15qqC67OuPTzbhAAlkyWZ57DBxcjshy66s53Oee8NfUdePW+qIM/rOU9RVqNMBxgGmJ0cJFN
BLtBkp7pJ4ts5AUrGLVbgC+bth8L7QuophYoSSYhK9LKwa7meE61c91AWR+GHlHJE4IHMONy83Xk
gN8fC4ED8GWm7/ksrPsxZEIK9VE94ItP+PVzuHtPoNIMCqZTE+r4pyNnqEVOY/x6SQj63Glm8sMQ
FMsqkKP6n1sWN2r3KrRsbqRdTB8Fkbmp/qRbDZsg24GQ45AdWLOKDScswu9DOeAaxVu/FGEG6vVP
1dLEqgKjhRUdVE9Q0ZwjZk0kq5ZmfKoCdKCmlcBZt1dLevKJu37TQBqNJW2SK6WkPt4O0L0yT+Eb
yQenXMV3d/QEJXapaIZ8Reg8f40aRhkn3eSug9w3sesTsAi+uNBlULt7uazortI8oi4L24K7unrF
xIaCwxlFk0xbmwIsnILL3xuKphDMqVyBoUk5zHJDZ8hT3KHFO+1De+RCVTd21U35Z24q1Ced5aLa
QuMOK/d4HytTSXY69f2IiOsZa2C7Vz25RgMCOuDMc5s+Pbkqpci6CWVzN7PDkpkw+K58gbO5mQbP
Pv4Tqv7fXV3uWfCssVq0uhfo6Rp1KAXiVy+hBR8fPCCX54vDQ9rbm3KxDcgGs6QJshnVqCynFW1B
93dFpOqnEQKB78uwnu3fdULjaF0uDhrvUmN0/N6X/CR4oAOGvm503S1tInE6gPcIgJ4uqZnlqrla
mhBUFghR8P7Hsfkt8/Xq6QkskU1BvMaMzzZ23clDd1kldXOAcPyMk5ROUm/m84IDtOrXO1IWcaUT
0wkYsEks9himZtjKCK46VIITEqkx8bvNVgyyXjp7cMZ87hpa7drJI0ZqYk4jRGcSD0+uwGyL2dAi
LRz7437ec+FUPIsB5sy8Hh/oLmK00Z5d/8UnTtZeG1Q06Q7oPb09ARRkQSKqNxbzdMrxrDeUEd7M
AzZRQCfmHun+EZaQQHnU1t5ZyEo+BPqiC6M+UEtRxc/J7q83hDbGJTfvGR1+fPA4FiQbzgcYemxS
9OYT/LpK1Eu3GNgGOAbb8tkT0+lBpC7gwR2MeREISlst+NlBUOa0ALxpXlx6YqI65GEGhDSxgdMO
DZ8ZDtvnEqvyLF3/xaZcgPmFtSjXsW67QC2BKjFDY+2kpx2/m5Zy8tzz/KFq8ONz/VR1W+4RAlWA
kkQh/YOlhjfgWtn2Sk+kH0IXiMZrTzNhTmYMP5bsD7y8JgU4IEJWr2JXeJ+CC3tXC9ztNCjFWIw4
Uk/56GWshxc4tsjy77k9ExoId1NTLo8J5rr2amVrWiRbWVi6FxIKKq6t404YGqgMtNW4oWvC+YQk
qzJ1kj+OvTRND0Py07YxLphIYBJIhU8NP0BrE/+qQb8f5npDUbP63eZZqsQ9LkCqnNbmz/7aQeQu
RMyim7GIRjK+aWrUv7oonldv7b4KR6WnhPC2ia0xWuAKNUKnQPdZVzWHQ67gOhZzkxfqoMrC89Vw
4jlt9sDfEyN6/dE3x8KiC6UMW/tpZO4Bw0/E7f417kQCX72rFVujRPQGN43wM7zc862VruYyCcUI
39rEZFbcXLPmzrIic+FfcqwfkowdMnV+YYQpTrmmtIJVLahUVSDD2L79vZGbhowNYa4OA6VICsQr
SL7SB6vvfV6FGXEI8E8J2xQQ2fL0KQidnFw53WPIsHhPMFvC8QLQEmT8A8NL3C1kEEmgzv2QXxWX
Yo2ulw69DWrAGIPDztOXQ4jZNlEgBO+3EEU3JCM0rz80v0H9EhMY5lNVVU5U/bIhlJtaIfDGmfFt
EErUfajVGJiWoOQBMkR+DuYjfSqRl10BmTuApvVAVpdY5V09FRg1j1udyMd3GFPgeZeBwE0YxHjy
mu+R9uv+hpIGi1/ue188xxQP5MtJI6KaZt9y2lAZqCpSFm+ousge/7AjC7nCUCTtxuj9mAFPfen2
ZkfRf9JckuKh7SY8ZkvkG3tePCQs3NQRAnaoSi9Arzu1G8AGCfvPthgHiyDsJntnvJ7BT8IZ+asK
5BwrBOATvZjCf8tZeiaeddYwvWfbLGiIEgP4qhgLGChOIynwisokMpxhDiNFpiSrCgrNnfjWIf5d
l9ZrWeSFE20mUFLkPWeELiz0Ha66lmnWQMe2qdb7QmDXYGwUOxTbsptkoutaQIR4W/Szf4jc0kwY
neShlT1EV3k/3qtbcYJA/7W5zH1bp/S4i66DtZln3avrDDRp54gMJpB3CwtF6Ox0TsXvVTCPTH/o
MnvFQC9eShB4daxsJfVHWQPvbNcF+qh44I4syepFyRjquGUu+QVJwWNxK2c4qpVgY0viwBEKyrcB
0jKDK+Si6Eso5avKI4MK0Y3dKsOanmfmM/p2wCf9TBl9OsrKMK2AACf1GQs4f1Yq8iWqE0qi8bqZ
xScDb1atxGmCnKzlqaOW0jHqisq01YMXSvorbfsPiJzM8zac99FAR579U2DGrbWMX4atCo9vNcYB
nGZGUPxUQCFZAbwdrzqGGladu/e9s9d93hqBcF28pGwFTeA8HTNS/vUA81hbgpkB09m+4QETmOmd
h2MQ9l5laaXyBnpuS0UG+dwcs+rNj2Pg5AnZc95hmWth/RnH8+c+izE8XFUA4woyBq3MEsVifQyK
ozsKYAsJ5acY7B7aW9SAE2HPPs1Uq+jkjS9/mKsTIFGZEw+kkemUD+XVttQ8sbbE6y9XrIIMRRf9
ijKrM6cpkRMVwHONBIPRt03JN8xkPLASVKLnJjYduCXfh4n5EQ+ZmUsE8mMeprWTcPTGCpuo6dUs
ZM7S1yZiSTBo0UQ5U0SORXYRHsz/4T2EoTborFlH7gfGS+fH+a0L5HxIRAckZtrIAOYEmR6dqd4d
vIsYRSlnkQJ44oDlvP1EdMhpA1nZT3675iv9JDnpvayw/0yEoiEIMhwPRxMFPEWl6NOmrzatS7XA
qhc2RZj0KR9P3az8fL20yWUPadrl47W4Ii3MrrLDSJxKx7ijcZa6FneSjnGiV2gc2wI9MwuUMWFm
YqHYPaoQXE67FYeIOOQdAJVxqwcBjmkkM99mb8fFXk01wxkWJwmQh1idVwOkPzohUkhAUGbSa73Z
KlNUCDOK303mw95oasgjMfUV1x+AV/5y0qkSo6fkCLuofe3ecZPiMDgBbd4pEcLP97iL6sIXYSeQ
sPHfp0cvJzgFydf6jIwzxzrNC4C1U9qPn+zdkjGTbL42j9oE8N5oW4Ik2aBZIge1vAL71anOJ55Z
2GiluJSJ/vadDWLlEQFNB1REwAKKePPru3lwdo7LlEps9JkVE1tdgQjHLvC96/OisnQYLC0ffsz1
auzpiHb/PywhgGHyVnSC3oz1RUVaF/1yCXe9Z3PlPW8McPo99pbzfASh4+eh9NtGfGYmMzEKCqtl
D1Jgmj8be3/00dpRRQIc7wARQEM0tOAFceGJgHkXXvXYNkng2Yqdsb530G42ci6f2w0SPyPzKFOc
PlNt76Cbmv+ETXAw0In9R8Ja8krElLuLayrA5J9P2Rhy2pY+jSCnZQYlvvxVzY9JVVZ7QP9XbuJa
X/nEAY0kdKvdvF3Vjpeo0fCMcyWKIHpeoTPg0EP5RSNnN/5rcVeMzMLJ/Cf2AKvsVLrQUAJVur7X
K2K8nnrB5qodkZ4csfvqyoz7rY43CjMPoa/A2Y4/dzerQXSjcuDn1SsL4ZO2B9LhmH+EyP9Vtfkc
zdLJc0CxYN3Y9BGnU8pXnbxmvXEYOq+cbUcMgqy60DHESNyZSnrfnCQx9M/OyJifzbVR1ffBYel/
YpBfc+54t7Pir2y1qJTcfc1fS0/hvQessqixa+HxwAFcUvvKhZEVzYuAdaT7gau3fqu4QMq0Fh2u
I2lAh0Y08o1g/VxwlukKSfDw7owO6+o76QO9yCZmphCUTC3TcOynvFbY/Pv19a4/MxQ3XA83gOHx
aNKYnR5Wu9dmRVABz44L+Sv9Xr5ng27nNCnG/g8VXYZASSyojaHouFSUHaH+MH8owMSQ1Q7PAVi5
o5aos+3XJ+q04TN0EZZbRCOVDLV4gVmXLEJwGTU/DvuXLbzipo5cUCXplJdyaCOGrcqI2V7vO9+j
DFn4u7/dAXzr6eoPxuoYuzynfr7iPgXNh/V4b1fDDtdMHu9e1EacmjOMHycLvgwrJ5fCSEviy2e6
bV7Q6aoZUUYRa9iqxwVz5A2fWVXfzvu8Mc/P63u6CDCSRwgJ+6Dt6UCqd6trfKmdK80yM8xKkcVq
N/7VeshFrsmjmg3Q5Vu6iHJwcZ+eLmzmDpqJtDZbyvsur/hsMrHd9hVq2x7212LKaxLVdFUmJFZW
MhaVq3L3aB9dhyABf2rd3evR/iWW4ShR5J2z1AhlZcNzzyaZ8z/74flMRPXEH3JbjkxqvK6scZH5
LDEstFVfIX9dFcqkGaF0BXEA4cveYNB3nn/dCpYfaPYs7KeJQoLV8EMfOHnQziN3frRmPuxbNAJm
Xi/2j6oUJA3c2ZNV5lABm6TXQuCgP//i1ay5a0y9JJxqFOtJHtEx7o/ciX+w7bMLI/UuIvjDWLBE
fE3jrGmJ7D6cmcg+49ST8RhhN9BT8Nxuq+9IRf7iocqbkI4hOftLIcKuql3yDHVykyWiCGW9dEgu
7zlJzgKJ6x12hSMbJ4+URFrsu6xExWBr7F/K61HglfTCu/JW3kfD2YnA/79ivK9oSHPmZSPZEV7p
XBixiEfQsx53btBMpasIKCvxO1HpIzZvj5oR06AVFcpDXWfykvYH/4w3uAkrd57pPpVqwcStb8z+
f/BPo4FUUiKChea7ZBEUFvMpwGl9RzNYsfFQ52AxWcCQNOv/ICOIAaSJ3uZHThILYzuAq49MLpUL
E3RcnaipT/1RWjRhdHSkIBi0RRgBUtC/p0eYSpoNn/ClNAsUqy3HFByBOwykM1p1VZs6E8V7uMla
DGhaRSSKeryJaAcfZThiPv2LSumDMubWPjoUi3e6VQJ7KuXO3lep1+LHz1oEUcFGpWyAvqyhFFqh
QfHlx5cNWhPDkbtHJVk2WqaNvZNVzH+UZsTPN+cZOvnzC0cjK6LawJDF6xUJ/xFW8WF2vU9by3+9
Tlt6rvNrRGuYuktzXVbZsMzD8mx41Ycjc/hsQAUQhm9RwBDXk1bdna4XhhTkse13ZV8TqnCdByjL
+Os+tn0ZhOFDs4Jje5dxKP3ottNBoJSj79L290FEyOcsISAZdU76VeLSuo5DL0fKi2WZq6mVO3mY
7PSXCw4r0FiN4SaozI0LuocG17ER8Cek5L5Ok33fXWde1mKBhnLxRnO8KLC9KphYZhn5bxVNEmCW
PRymEV3Ocpx5CwKOqpQ8c8JOLpyZHc6fniafTlgBwB06jic3X75U5QmEvLb2jZm+RPUJLOe8FHJG
VjDri3SYufJtlLm+nZraKru6RJSUWx16DgM1SYc/0YKkpwwySsml2SQfLGrzS/JZBf3uHMJS8FLP
5vkyTfwNF2/dvM42w2udcZHbpIjncIbMUQiHRuBPnhI4qKDPYm1a0WaYgaYSRyUqWUiqoi/JkUvt
EJsVHPF0ltpBlpBBpisMAk9T/gTfEb+xg47uV9YNin/LVow60ruOCQuL6WYs6RzGFF/1Pox7Lp1c
wes6mZ3lj+rRiBbP4KDT9bT1SYg3+VCVDNpEj8KJzipGJzbDgYK68MsS7bWXYDOtuJGSB0qRifAv
EkFqf46oyVY6kGkZHeUms6+xXjvD6u6Avfo5Fn4Cc6wFJz5eR/3vpmcElXrEW9pTNADLxonq8jjg
9OMmNTJqF4NAdCXv0+WZPC04XoUTx38JEyccJvsoxBh3u0NZLYSaVR+bOfxVF4/SUX7R4nHBq9Tz
ipUO7zapY5zrCVjbot1lzuXaBiKQyNocyO/sa6rdEsPAH6C0axJ/wavR98xVuSwwqJfO9LZGULOr
Zxv50ExYliUUtAWe0unBrqzKIWybVjG9Q6N/m63IOM5zTKTRR0kir0seSpBzz7E4XSyiqLPKF49R
37ShOxQdnN5JbA1x6xSTJ8T01p3pMSsPPmgmXQH1vCGM5OJofFMWjmN6UwQ8Uer64EEHRB/YOrlm
W5pOCHd66MCX7weqPCm19DicYvH93Z8YUNUnn5kF6RZmNDDoXw26sorZD6+PEdJkjcM5psknf4yL
nWYEKsYVRvKXcm1Qj3QCXFy7K9n60fHtTuttmOMnoBPYIrcBCHPGR7rYyPDqwOGs8sg2VDT09LQB
qxmJVC8nER6q1VlAE3cgwQ26YNtn09KDkYpZjeQxNXmRIK7kiqwzSBsxvG/Tq1JXGPR59g6k0ISz
OrTKRwhtYP89CO97IltInTSf5OEtlLMaAl1UKiCHSR2oIJtuzduTJsOadEgdvmfd5C7Ye25QYkW1
7ChSYC+Lb2Do7edC/G3Nnf8EFTNsE7exytuRwouQVFuNZiWXAHojCawI6bwMtO/e4un9jZZuzzl0
vs5aPslxI1AmzXNOP/Iy0RJ55lXyAYf+TtwEmGUFJnSVJLXnkDuQmjCpY9Cys/XfRrfHQ5VJOMUA
p7rOPxD3CbnCjcyvXSfcvMLnoY5riGwBFIMaxDdW4MlmAtn7Eh/Gz0DRMHee4+ZkMjzrVQF7emzR
8cxrAIqzG9neGQJ8abO/7GSazlSywiHElVKDB2ub1wP9k/L5+7S7s04XeUJ6bJpQ7/YiDs072/yg
BQeUmextNVwmhLjTwKKf01ibsiX8oCtVkhhoeobt9fdxWQiLwCwkC3mrxeOEV5SU+6Xv8d2sBTos
jDz1VPbvV0X2NMcDh3h4vFEojjwj3V+ghC0P5r/lOC5tKGHj/W1kNmyIU08EJcqfDf0TyW14wgXx
qBKP+r4Q1pPcf3QLcN5Oupq+OIk0wWk7ggD6IH4LHlXwhKPerYieoT0SKgOYe+1O+kfgCtXgziaA
Anz0Ivw+cbgiL7jC9ai6SwHDVA210u/BCZqcKkbtyhsa1Qsej8alShFF5pBmeUoM3divo2c3X/zN
yoxpPikGnuvGQV9N6CblIgn+j383oGHIF3fl6kJFHCL0UnYGL6ZKbrZxVNUcFLAuSYserrc6bTlR
Hu9meqtjTaDWLlJGnSkpMbNwkmxDHKDe4IGm+SlfpgZ9Xeu5DdtEv02rp+ylI9nqE+LytKmC9S4E
ey71QbWZt/pltfiODs3ygEnrIjxF9FXwJ34oj7jAu7U7CWJYu5K67O9E/JFVqCdLyqsMduHIDhNM
j80hoNLQtdW01OIlebwbR7mE2203Qb4JHOxbRFfpwENfBwypwn5LXEVVKqFtXxtaVJY8B2gsKfab
xSuZ4majWTRDri4XpY3f8hLRijwOF5lFXDe8Cny3/ApQJYo2GVkeD9HFpSuO7j8EZ/MENq//iTx0
pHGZQbxw9gg7yg7jUr51BdJd76oPt1kvRJHUDjkfsUvcEVkVi2YSUas92RwKRXFhVwynjSJ2ah+d
7ccSxtP8cUAt9MNK92PjzhIm2Q4o42II5mLhJyxtcrP5Jj8htVbonuOgVxLUcRv1rI5VZmzAL3/z
YrGZc8pjEVwJlQ2VZBDcB9rOR2/F/cJKNcFGaiqMnO58fqNm+SiA3KaBFV96otIIqofPTnWu1ir6
s3M3LbcoUdBB7vbiQ3rFs0RfJOAnJ1NucJzPjUSimofhGLgZIVbX07Apoz0+u0bABsDI1TPa0Zcs
K9T6oPexsXnOHD7/09YMMha6A1TCX2uT3wPACAdZbhPI6X1XpRv5kwALRPJtrz/pqg9Zmc8z65uL
Cy9H0pJNwzPfvB8Xa/9RyFiMi3EiRj65h+Nly/UPVninmdCN2jhYn7UQzBuhzB4d6Yq+x9zvj+H6
wsvnwzeAtKH9zrapwshzSTRXvX86KdWeTe2kYfcwcKvN7TsBznFzGyEV8LXVetLayUaqJaXAysh2
9l5wxqCnOtQNGULLvyG4Sq7Tq7cUeFKTTNZE9maIKE1YCmZVrxTNPRi9yHYy2YSFTFP6VmoomnU2
MgDb+9V9jrgK3erS+s+IKu5htwvo+HEjG5fvQ2ztci2/RhWXqdmZeWwVyCYC6cuGfwRpf5oXQy+L
eOiXp/4ZSpH5qi37AcAFtT2J9J+gZ0AQ9xiYTnlYHEZJvx5xd8h7CB/IIdgvu5ATemvc8DIvc9WH
r0btviiHRwDv4V9FiYtDEBUBRvwakQz8VE6Y1LYp+fZlzqvkixIjRWExEVwzvHcuMFWGOqcP3lsG
qZ5P5Pb9tUDNDaMuh2a31QXUHwPSrvqprxqbREmTxXQHt2os2pVb2rXTUyA5lzwX/Zzuk0yTqOij
hA9z/HRsWrq1M8gfWSXRLzTm2iPsTtXhUCmQemiE6j/Sd2N4FelHlIybccXkHY8Pjfjs06WIBVTV
bBjeGTO7bsS+zKBSkA5yYcVprFUiiEl/NdHm9z0QEt+7Kfyyl1Ei3AJDPifdR9xgTgSRcsczr2PE
FtO/OKW23CFliUjgnyEBNe7Z5TTjMo0wtxbNkhjcKsL0hCbonnuVaAT8REwNENIsGhELRXCCtzVm
K0CU6emfKu62FpU9DfV2sDwx0qrUbZTKE0m8GgEVH+89cXEu1OSXgD4ff8/NIAA1juyoBmRg/p/n
/vSGc79T2Emlumfijauv9jq8t+z7PAuoZyoMNZu9d0S6oIn8PKKDTMcWUqSsUn6lX9XYirSV4t4O
Hy5yFqwJoQBPIqkwBj+AtwqN7XZx9oS5ThiSxPXDewKSCtrMzlAEBF0NLIrKFdMCXrrjzpSuU2GT
sfjQQguv+F7QBc1Z8ennCbpeaWraqXwoBlKS0cDNAM8TZZ4jkiRUPt/bcK7/VTvpY1/qMcCdrXE2
VGG8Y8BdKHjiD+aAgRaZ5YKfoqs5BYljbKyvauw0A+nRFq0eOnK8+zXKKfczCTjlfXSxWeKgxMon
gL3UPklaEjM99GLO5lQW+k4C3BJcOWrW4ReYyWMHbATYRA1vPObCykLc7qOdp2YtRYrLgHn+A1ww
bW4zVfvxXd/HIJ1MqcY1uid+mfn2DnkR/Hjc6Jucjx4tBhHxtUTnesZhOwmCd4gv4EksGnDYQl0Q
fqt1bmdLcITtvAuIi1eE+Lag4kpRcJwsWIngrw16mXKCFq3lol81OLtrLVbBCbWIBa35OmDfbz47
fUKTrbjTfrmIq3Gtrnbe0UPR1p/9nE7T4ETUknjh3V2naMiAdE45gSY9e7UWyW/9FL2oqYi0juO8
u4mvzOA/d4FeOefuAoKRnPjuzibfTVE8S4KVUPogyU0jZc34JzQIuCjwW/nCY/jrdZsOOjSSHwEv
nHmezdbazynBmgzaUgsYVZqac0rHTenH54NGlXsMrmLvMp+41ZE0eA3fsCnwepBnlBUaxgapoFUe
vtcmtWN7fBNBZCJELP9zsPKmEEC9XWPetjGxocGqa3nrGZfdcsi2uDze+KTUn66AaGUfddTRSsJs
lT6FDCwPqdsqpMT/5rQ2AXoNjsWlwqOouXizb24/4B0RZi4u8/e9bAojVfaYYng6NaZaWXXIUYqr
KTPC42xTE7puXQTzlVIxDCDN25VzsSPWpDThQugcBN6Vbb17r/mh8ivUrPL2d+dIXVcJDlHw7KQq
fw6QtyUKYjeckDVFeXTuwIJbxaUdBIjIjxDPy4tF1nWWXR4l3PbYtPXTljWKb73aq37LH8B9uMsY
S0ad+9BwveO/TAtSgGbPqFCZ0pnJfArXHs779uaP0sR+eHCG2BeYYC29JKYI46xgX6we81WDdG3u
dCdbOO5kj1e/3PGzjYegkdkp9uj7v6HTWa1TDP3302g3QmAe/KWc8H8MGU1kooTppEulS8zhK37A
2sLEQJAmorVuVcIWc/4vJ2izXVvfENguCRS/mSunnjM+xdpxzwGL+C87wQLH1Efps6xuOMLP3+yA
eFZknICP24CHPgIgtMDhVXtfJev7Ltlnq0S7k0+EJGZ+QaEJ3c0GitEpn0Oym3/G3nghpPXN9k4Z
dCfGj+HN2WmlX10N7wioHCSkrZtd2+lmoaPniuUUyhD/fTI9fWgOFbYYT7XsImiXcyge/FvP58ZN
rXGjuSe083U5N9GK98ludT3gC7/GvZ22rf1n/Jn1dNXq6BMzhyqPINVo4nKSLXKsMLHgXdI1TpC8
PXvIA/WjcmYliiD0R+2DSbI2EA0tMB2pB/l9Pp8889xRJSjZwdArEv2JC9h2rRrHbXrQpTJaVM+n
B4eipgpzfGnrt/UgMhI8/sL6hhLsW62GnlV+NV+7cLcrINVVIyjAKhrT3QUMiDmxAThquugEcGIN
ggUiuRXGclQKeEyBdsilN5FI7ejFKiA6/yPq4KiwpfzUXq6jz+sPkFBdFHw/2Gqk7AeC/7fCPgQG
Y3Axiy3fMv4IWfyyJrTpRv5B4YD7/VqYOu4PBl3xkUs9xhftSXAygwUFDwMVU2qjVQB8hRDZ1Ar8
UdBt1DwH0KrFvjgucB9nLcKe9Yk5A2SghcfR93k7imneOa42lO2Vkmdylt5A4qOJZLs8AKoEJF/4
LE0w2uOq0O8pxOvlJnD/4qOQFfsJOdzLoOsscWomtHeG/1wBD09WM9wOcvYx3rvHXfled5Mjr+fz
hM6M11A7oASAnh5GUAyb6VG6qMS4ViZB4EeHfArFmw4IFzUMe3v7cckk2PgKiWO6ZFBLdgEQ72us
pQeM44nmfziqqWMsaYUtaGQqI2ozskWz1i5vwZv/nyrK1foU+hLuz6yIBqqdgzn6hmY9vZOLCIsZ
95kcNA7dvk8gVn8SWPMhD3eSHQckGfSpxx0ERnIWUqNGU0kwziWKV3gEgL4P0g2J5KuqdX+poKdV
ewyC+D4lZ7lsSMVVQFx6y3WuOUiZyG4EV8iVncLUJNZ6PEJS5mtNAylD/ccWRSpzuPv+61kEC1SI
iRWQHGD2OMoBqNWXhl2dGhCD5pAs5ogJk5JnUhTL+Xxqz5JcZbzEe26h3vBXN30LdrmrkMh4B1tg
/o4PMUAoK7d2Weez5yfmp1j5r9x3xDZJ702FKJ7u2S6LsIXJBs/JNuByCjI1WwCsK9bm656LbDj4
mItIe6o71PtLlevrHzI7KHlKelklfywnrBM3p6oaKwE6oGDbpUOPkzs3ezJMinr7/X79vu7GRW/W
I+C3js2e9Zm2blz68i/68ubAYiWBNK56H2P7XGGut0DM6uSe0a5gVFtcG/y/bRo9rBxezoWdNkXA
bvzEdWhOCjkuvbuE4bPvLsjOCTPOm4Ijs9hQtkfG2fkz8vHWeKErVOMQU4ZIfCmwbnYgMqENhmsW
LWhqU9+rSriMhkMEsB+7lDsgMoasfbfqh7bCpLLEuQS9ce47asCDFPmst14kLtpoDnhjg0elan7g
U4S9mP9eLcOgiPm4Mj5oKKzQzG9M1kMrxRmg64DHuChWRFHms8AXGi9OKZljQuu5/FtzHLc+Rjtr
jmaRy96/wWLG7uIiCwSmoeJiLDr8srIDvYBKhGG0IcFMxV/WmLEJYRU+Ciz7ERPaHO65HnY/Id7I
rhuJXCbxIQLRdNuSIly+njABkfnKLCVYZ52FAp7Mr9R5I321NchEiWoLUtkSBO2ek1MbztX+d9AC
6m642i0nbmBp3n246GtXgfgnUCooJ7p5FrNDLLUfZb8Ss9mcW1LY4Lc5PQiGKHUDHc1NWXLj2VgT
ugHa7tOW2PHFRQHN7dSeoClaxG8wTVonJf6J9Vvl/6vWURmb5lOubcpWllr5hoj/m+iU4NuoYD4Y
SrtglcKVyl9AkU584pfLJHoxBQ4td2XsCI6vVUfc93C/HrqCif2z5gIRcQ2rfRNSXzz/4CWC8JAr
j7Eyi37ctSZTj6KBpvJeFWNCqENZIcKS4yiZPSyD2f/w71a8shE0Ko5WPxxL4rHVFEtyIUTO+cWs
NF8MzBhMAPfzgXtVPzgWmDZuyG4eOLZD9iHES0ivFhnyPHXQr1He6vOEGHT2P2pm8B1ny8lbLFsY
mF19XrISHaF+HT/Ok/yrRTt1x471ONeCoVcXweyyPBYh7O99C3kH5ErW/Nn4kqISazmWiw7QzeqO
I/HkogVSZsV1cmBkfc67cgz/iXohIWNF/iUvJtZ1OrW7DuaS9dG+MKeWPuyhkAliwI5Ca0614k4w
2fzCaMgDGer3uplSKF+4YvTsqBsYVMpIX7V+L5Ez3VeXjLlpMPLyVkGyoSHUNgd9wNoAfN+5vwPj
KdecSEDFWTt88JHsb4k/xNwHlzcV/i3AMsF4VUB3LaNYevh6gmrsB9LLDCU8QDTHhWjSQYPolyGh
lpmqVA65VK/B07EByhLkruYr0LST110Z7SlFkA6dwLYywuKicOMXshkumUZ7zYu9RpY+bS8A1eGO
5ddKBLVZTrpjem+5kk1PTR+CHsfgOztRdTVomWyLNQrdKZlowVTIrplIUIFPrj0CBgTc3yNQ6YSj
jG7uN4ob5IP7cIzyuU3cy0Jh4mexjlyB4tiNSSiNn26ABEqcMjCxhwFLiADWtKmaXOgFBoT2PWLp
ETXJ8WLpvDsDqvB6V23edFmJfiZueCXsn0bkhjbhT1B4J5D16e9aVRkICdGt3rF6mH1JfgMNEFC0
xNk5Cy21quuUlbwDf1sobfiBsMrzYVNAVuAdMGbC9ZydLplbgdqPyNAJIL1m1Kb9WVLLHTCnAOIE
/fueERuViyAm5FyohMC5b5/qb2lSsM/pztDMi3iezwTDp/VPPgZrzGvTFKwHyncr2K9j94Pf2L+E
iwNWZ0bsKXNWIf4aWDoyh7v+rrjQn8iUfrmUwc9/EeGFt+SbGuWwafRHuQ62VR0it5c83yO4M0XQ
dJp1XaEbaSzVa5Yze8KLhgvFF5SuPthE9R9ntCRjZ2h2B7aUEoDAqtVhpzmaRq+b8xsiQTHsm69T
6IFPj8gbAgzK9XWkXfxif2Jm6wzS8mvrgAa3rzZljE//8Q1BRMQ5h6iayhbcDF5lSdiSHE6dy5nW
ThWaFsn5SHK7T6oBIuQaZoikUxJn1az5b0G6r7TKurGOBGnNbGTmCl2uRyhTcNn/RFzKTqbACJ00
nLHhMSrrzKmwnAiRYyb7mQylhMmxJw+nWUITljH7pyd2KBkkgEMkaYMLSebf28NXnpz2rLObDHMR
12VpEtloTS/djx+XCIjiLklhkpNiUKMr8cSSmxGDWo/+IK05YaicEkwbUwViZrskZTh6xTUYgzyk
r1AYGb03aAe9P5F+en5PWDuH0jQOhtzXNvzXvrqVVLGAO5L2/7MIDqUYclcvwwow5qgqf2KWnWvB
+5dLC6RgS7SAuN8Sj7rtJdr3PGqNkI6we2kr/1vucVpa9SHhrqOIVRQbal7LCKQ+e0IE3FBmxjhD
bcWneTsIJVMWzpGMfiQslXYQffuEZt5AjrqEL7tGLjxzwLc71kJooOTsWqpsqhGovu5LAqQXFaAY
ntqxTOb7ygERnhpgNisAV2B5d+pP+PhF+E1Cg/y+XecAi8IjFW+OcpK2rLzmSnK205YgIzUXrLQb
0iqiIWYJzxZdsCsx1kSgWSArlPvwcZyR+TivVLMsluJhw3ccSXCLhnib+VvtvpMUzTUgiqGoE9i/
UGwvopTcuDVL8TPn4+7pjlWb7P0Ycr4uYpY0z3v9TWfN1DFXWB69SZ1+wbLlz1l6UkXgs7YCDdq+
fen4eNlYkgVzA8hu7YWUouD4q63d+7pd66g08mKitEsJlD1MBvOVSCBGnxXAh36JWR4jvFXLoZ+b
Dc8WiGHsHYHdPI8q3POpmklPgkviIodWThlEnPh4qZ6nn2NIDdLfr01diuFuSNBeAwtuFAtpEP6K
hXjqEgklY0AMk3ypCzpaB1NraHz0WtZdg6YXi+3X4IbKMh3t0fX82Bg6ZdyULq6V/PGRj0BOekXn
uZ0AQRKwUBXAJfQgTkB3ItbsIV1YYS/PN8inuc87Vi/3L2oPiS8rt0nH3d5KMM/rZtOstYi0Poe3
PQRneE9JFsvgtyoXvSNeLdISzdklOmIFwQ2tL729m+/sbKMyxGuaEDVQs1pUolh5GyZZibje61XS
/cjnHe0zRlqi6LXP7oqvDwj4TDrvxcOTFKaeVPKcTqLpWai8R2r8ljCyO0tKkI5ryc6kixSWte94
MihcPqmjk9S1yzhVqcI+bY+4ROe6kq3UzXyjpNSBN91KvxnP1BcRiiFP4uvBxYSgH96B7/D8Ukt7
GK5HZS5VUhNahkoHHC8AkF08z2BZEM7Zyytru48ApK4Szymgk9GN+y9FOlN3czWwWnLOSv8je7KU
3Icy/V5Ne5mLRJr8fNkwl0OykDg5KFalmNdxNRjrqDrFn1P43YdHw4jFOG0uJ0RPEuxSmiX7azYQ
ZxRSH/3Em3AaO5Zh75PADFLqliYQSgPKhbDlB2FyIzCBCvEVJnGa1SMi/9JgTnRsJfwbwa9KjeG3
t7ggBHWGEfhAV1SSBrNk2Ig77jy91DRPy9Vx+mpa3psGlpwi90FcQril3nZ2f1qCxJW2Pw1SJfCZ
pjL+f+VnMnEit2YhP5u5ArCMBsgjYTrKX3V1Vd0yqSanbE3Iq2VqFEb0c415pwE+WcSOg8igI9uB
7ZmAbnw4wd2+y7eCACjbOCcSVYbxnWp1t5TAZ2Ne/heH6poawG21gqA2Qq8O3KrJdDF/JaSYlLvl
gdTOXI4QIsJyrDVrzmyzGc1P2zq4wbj2uz0eTARLddjnKRTna/1KSjzoUPMd+j0r6N4/UoqQbA9U
Vp9ZXCO+vhDuEIj2BoEixirQDI153mBTjFy+taCezQ/I1siiQesYo0R04uA8nn1qlKG5w7DzKJey
Xb0xLqEJug9aesZshTAxFS4IVGZjFWli1F0CD+SYwsrnMDhYejCkWFOKgrivUKmlVqG2Yd4Y3ZJZ
ccSjgu6bY0TuJMMkbdFJmgkv3i8IVzcTwYjOY6MIi2WgCwNbRXfA5MHoJaIlQTWSIqD9gmKKBRQb
0kntU0S9zQ0+Jh9jYAKmQp5JpSjplqWzP4tv0+2VHk0hM8QmtCCP4zRVKwERJJK5KAiq6X8A8iRw
dE7M8xmBER1G8FGUDAmT73Nd0kZ7K7LtS1jJ8N2xL9ivDxDiYlCVlHBZ2+2pEdLpo2EQnDAoIVb4
jFLq5NzdVvdOuVAj+nJhOV8NStXn4GXZHqQJBOhkvoBoonBuOv9Pp1hiNP2KiJwDut37eRDen4ll
uwB5QlUtd1464iyBCSG0AV26cxQUmWc9dHbjkM34SRaVG5769Pk0bPFmo6esSEQ01GXA8hMK1RZ8
UOSFfWzJ+WYFLy4u2DaXMld/fa/UHFj3wU7JUIqAbpwA4htJFZFv6v7jSk3LcfP3OtOpMuNEeS3Q
kBNCVEUa8Xo1e5t/Me2TRztvbzx+rHaJVXyLbFQ2PRn/T/vxx1FGObg4HBZNsr6O3N0deivKUXkw
4apgxWjWSpD6fapmo8zwDrUfFi8kctrq2zZiUtW39N5Ui5nUC50pjz9kXtCdsNMb59dbPIuxsmOk
biY8M8gUYCmShKW2F9/Qz6yR4wVjvWphi20+vzMKUi13GELmzewwb1J7NBFUFxo30aIQShc20L7N
GXItZKyWn5v/cTCWjTODYQ5ndz7FwfSOy43qH/SZ2Xtb1BIXNBr2NuAgMH45cYcSxarAZDlBapck
iCmhvpReOpM2ZYU9uE0C19ebZb4nJ7P+V6VOAL2RGHPP3FCMEzmLjEvikXCCI0LBYVVnBf40cuVG
OtuTqHWbop/qYHGBze9ZIfy6Ztgjotulo1WAdrmWGBhZvHmJBWkz7gtT3VvJb5vdJkWwPKqD0I9X
KHEa5NzAkPQgYAHg7Dn+kTnziZPbaTKCeX93BUJ4Am5wi6gpISsHqCWp1CArZBqmdwcPfs7lyIsm
zrdv+LbLfg9jRjbDxTHVYrXKbaOE3DPLPvHGcUhbGV3knpkQrZuelG5sk4j44uv/3X5vT0T7s0Jb
oW5HCxpeb+QpK6sLPrTvqjPMDm2itqeRJE3mbwOvXT2pOssFbz4x2YejNKP93GC0/tKy9bCkYlJe
yt8HuIbu0Ua6RdeHbjxa70/4bNIdUII22hibJmdd5hOBZdwQ7SOdwGhbZA7knwh5dTfpOuj7987y
P1bukV53Qj0N5eEtMljC39XBxXs0fhRpIwmzP46AyCCIGDtXGuluA4yaFqiGGsZt8PiqoHdTl861
gM/GHphb/JPdHZA14G5wycoNF3RR2svMpW2bq8v1TYHI+hltMAR0LKWCw1mAMcNlFoRW3C6OoFtP
aq6/aSsBNm+tMApQu75KCC8r3C6RbpYeXUQMtzyNXcl38rCHNqBfb1QmxxV0ArmPY/kHWhC3yWgx
E8KXc1ZIbkmH6/f2GK/9JZ6Kg4dcevxAN+UAfmvPUZUTm2qQXXJQM0cCSNTtDPPBAZND2yCHdr+r
11xqHbyx/aixaNPgSkVf6CTbfnLl9qhYtTjUhrTnaoZGB97/amlIrT9JlpI7DjUGvn9ADg3WXHF3
X3BWMW4Oy8jyZWp/hVI4rKxNI5OQC7SWpb796KW27dXisw8ypoC/EaKpht6kM614Rpx27MYGwnnT
uf6fegl/9hlGIaZO1ZaScKOkBFVKaAIJpjZ0jZ13ZMGgobBXkJVXYS2oKZ1zvu585O3YFk6BabdC
WnGdrKHObxYXFf96aGecQiROPSLVhfW5BWqAx2UGGFcyOhPYsVQToNdf1pGPHmljsD7bLmEDScTX
N8oi8kl7j5NvKLtvLf99yhAl/rTE3YXGZVC1HjcogKb5Ffwfcd9SU9VGUJ04kVtxw5OzFpZGgvOS
8WLHJa4vpllbPSD0M6DJc9mrjtiiFZ9z+CvtjW3m//BfC45/rUjIliBnKtlD/gX8wNqApyA09BpX
akdE/yjI5UTH0wXKCpXbrHLBV4OnoJJ/YbZt9sf3TClHCCSvCXRVLLYHijX7Aj3LK10vDSFfPcGw
WtJUOGsccbrVgQ9XFBNxOFzaXvv1dYhTJJwJteS2c7KcwQ75LCsUETebql+5RcYMHUCwXzDpIa38
XaibBaSPBBrc67H3kiL69qyrDuu/biByH4fnjWuyXq/iiGWun31Z15bVHG7HzAh856uJwGSiHYgh
c1qQ1xc8hgCCqiCbNcY/IFS4/kC/rOj3GPMJl22FeYqLWpE48rgKpZFquaNuChIGk9r3oEPpY0Fh
h6SMJodkcgVZK4QeeqG57b6+m9Evetp9NEF5hljq+YZrRDEqMwbN2OFXUpUEA6gRtAM9mrOAFOmI
WPEVcOXyRyUyVSzxZ/e2FM4OjKaIlW12rV6F7RwE/CIGXOwNSTko9pt7QU0JfUio0xv8p5BrxH+E
7uC+TvZoa8PBis6nAW3yGURo1Xkb79SqmEcPkK8AWqChHzuxYXYIoPDIEkQvlZ/XdtX3B++q239b
KQ6wPYarMFagRoE38Vt3ON75Z0uqUH/LQVaKj2W9DD2Zb2lgZt0NnynHw+q5MxtkwhW4p7UC6sJU
vc9Yjw5H5vI6nD2znvbhr+iMtYPn8P3B46hJXROyIJjG4UwryoW47RRxaU6mdZ5XKBJ7/9k5tsjM
ORpoatJWSpNxdrXOxt2EkfGXGrmQZ5ecWbvugq2ytYf6W7s4ak69UCZxg64hTJCnPrErzQRcr629
RwWf92kujN6toF5NjyvUXyvgktlV6qHDLsi+IbSomtXUGbPAgo8wfyjoX3G4sFRGUcoY2rCqtXdy
r6CdiQ4rFMVzUXbP/QA5zFxkLOWzhmOihCe4vnHyS0aorGlG+eZsKNqnMsR7mhbPjiMAFQqzZbM9
BI3/3Uvvw9tfJXi34bUAKOKDRchceaEvoZ+a1YwIXZu6xlqi+J/zvdjoOy/xmHiwVZu9TjtubFJ+
pVnKQbEPgXnjI0y1f5EySMT2RI4AfyZLOPnX8rtnHmMl1XwMiklQO+LYu4S2G5AEnY12SBuvNI2n
cpqS/R2XVqNIdbGTIN/QNr303Mth5iLL9OkSB5RHdthsdt4AL6bfAkKBCG3dVNP0c4RqTv0HyGfh
q85yqoe+U2faK/q4JahYE9LQfarQR1LW+7yftPTqMQ5ZeO2QdHou4qAs5VNP0ipNpjSSItlvy+Vh
vWHLxbChFlTNUnSN5QQnNhhc1hzbK5W3wrZs2kT7xi1LdigCeYhOJ6mcvYrIi55Hl4AszT1hkPuh
danjcFtrNv5VoUlBAIg6QMkANyayBamCUXEOfvMV3nJmC3kOGdwaylSzRhZGqGD1OAILvHcPPA2m
uWNVVQQj8XPN8Iq6erJ04R7Gu5JsbZcJJbmzCSZ9U5kDxtMlFAjM2OELu8BKDA6ln+lo4GG6lK0k
TrnmfGlRnKIY3Z7ulFC1k9iQMwJDqs1Lg4YxRpgeZAOGSeuzvA3/TWOLpWlulCpk5Wd7KtOc0/BV
FraVZlhkzIDBZpXUtkyVCcUoLWlTxWx+qpZC/WVKEpg0pWv9F9LcR8NvVTkfy+xOOMfe3cZIHp6E
MUoqekZmNkD35Qmt3aVPir4QIhejA20RQCbJDiFK0RfnybvWLCP1k1xwMSIVqJqRnSq4ZhM3KyFl
iyvuEJ+G9K4gKQwZGl5t/B4Huq0aVskHdQkUYRtB9KMfauVY20LPPU0/49caFgO2hvzG6+iwz/zW
+q2bv4lINSOJNfAkCYNm50a2PLoFYGkZV9+JIUoVcjCWLRaFLcN0zNmBDfE/+W2H88qh+KM63jLL
X4d2pa2T2F7CrsFaXmN3SqWeI5XlKE+QRvQpoVg9RJTr1YBKVdzK6JjeavP8QvaWPWjDfvW/jn+4
tM+CbkTrtAsIbDm/odb8CJs035wLkM4rtWc9fg6OaCR1+zTIVfaFWOyVExNgBgRWvGsfh4GQf/tF
qvRfMkLYsA5LkGC62hv2Xk0EnGmbafXKTcBlTlX/tg7OsbE0TAA8CKY7swKKsxQOAkYVLUvDeME/
utc6QsVEMCAzHN3+tVbDTXAeOaQFBJPOsi6OmREYfZTdi7kmRQnRKiu9BudpyERUZr8FkoxI8doc
TxzQvXTwO0d0P3tLKtSJCm0XNcF9Uhihhi0d+xMGiPQqTMo1Q9iV4sN+jxd1sXlP59uz8fOCXanl
IB2OQ1Swax5gRb+0A9GGliZd+6gOes9I4aU3XrNQEI2TqTWwRw5Pgb6JRaVl7yOMTzPM9JptkUzg
eichRWPN8PGN4nmVt4lmd6l25O+KXyBszBn/eDEH3OsJLFxOswQ3H2pkcYJrhKJNFzMokNDIZzQj
POaM4JM28J3wu2rZgDhPZGXf+blXHCA/ynvdCeaiNgGYOhicCcyzBQJYcCNzjyf4F0bMIXxPspmy
aqYnthsGGadfLlpiPwbHlFEkxqxrxeZ3/MD1Axbve1Vc65nB/HsLN3tPDaAWzQjd4O9akQCHmOPS
Aa+Gvto6vAki/MvqdhhmeZh5Jlcw3PiBCS4WgJ44F0EwyD7/FyKkHtTbbLJK0SwsqvFHxsQo2kTM
H3Xhl+E82GQmfIigCK/wrzNRLjAMphAIhkSvOl440KDha0TDQWiTM4BLU7aipuLplO3icx+yRDqd
IdGWBw8/pDCrqz2W6KAkC5S7tp7l+uG2uoXHtGFTMQSlKQK2Zgufr/9ziIveNGqlSj3fweEs7QHM
Kv/OVV1w5xpjz35gdyosPoG657IdQkfHJeIGKxe3MOarVvCcvOvbNH7kiuVibg00erwZovTPwWYz
v5BLc5wOCH9CBRhYnR2vKRhegLfb5TPNakBaeydad+GhVowCYXOSNJI0Bo9b3YjFWODbxciHEvIK
gZeVnOI9lK+yRBcKKbadAsswzrcE898mgRtmlR2Y240Byn0nAUexrED7la73zqU5mwutX+gRtP47
GOg8KG8A05bTGyRvm2Owr/tbShVbdGUmlrfswISjlQtpiEmyV2ORH29uxrCk2YcQvCBO/pApf8la
ZJy+9tEeodS4CTlJKxE/2IOxbLsjDaX+9K0Q87qi8wEdcMxb430nM3dXoLErnYHqdMmNdo7oFpNi
ieJEZNV+MttDK2JimU5g9KuegNPPzeMdfuZiOegoCZLMgwYvyji+lbT2WDRz62aWmZzmP10ZnW4K
wbZ+Vppmud8oyzlDR2n80IO3TCrltUh2R3aMm8yqZF/X35Mfc0ymvuJraph4IAlFPwUpDKvdtFSa
azkl+AY3aYyuQcmS0CmJRb7vaxRiPhM/yZPgnls5l5lB7dDWPb9OyILPs9I8mlOpUPSu+dEjbHc+
gOM0TvDpkbMMKDShRx+LR8P5GaSLwVorUxXYmmYjijDHMOEA0qyR39xsSAKq/NOGpGjEHxF0v9fH
lDqB4hNgoMafJ87p7pKLshVUtVEXjV9ohQX9TNeyLSHtUlde8JlsYX7xlZ7sFQMvCzLt6sEJlKBo
DoBkcCEH6+H6ZVUUsqRhFw5+hgtaaz2R2MBUdxmtvt9pi80nCoDU1VSfulNZrScNKQB3BU3g8Q7s
RM7sOWvVTn0MLldzl836wpEhS2QpmwQ3JdeXV8iWT7UH079V7aKIa2mclWaKCd+umM6AXOVWPXIA
Gas9/BSRSSzvbwbcgaqWCDDCOiMwSdTX0ziUdO+ocrfavfvSzxsaCzmX9oBwfyekX7wT0l/ojDPC
sUvOHdmgwRXstuaNFqPwbKfmb1OYfoPYGEN23WuziSWuPB1KqvRxg8YOk6vk/svMOERMMJwKRwhz
gOuoOjZUrl8BpqFxXFq+8nymA6WgYjAlCd64ZVOAcQpi3cherI6hSXUhW1is3j6nfjaFldgt5Y7F
6e7wpOoyZ0Uwpqkqdp/7owmWy2GZRLSL6AsccyJGaftzjzrsiNj5qcG6iNZ3LYlY9Mq9W33rh9M9
pvavP6uUN4hMYTCUuUG9q4anYO+VwJrrawlCmCVXGh09HW2JpQ9JaqRBt4RimAIQ8oY9n3qH+Mna
E2X/6u/H9YNWEgWg60l+AVIZAYh7NG2tmOrwpyO6606Ob5nb629OcqRzfAmYJh9vf/9Iyc8fK3pv
56GmLHvFQ1bD3Q+s7qfh4nmL6XLnHmb250ve9zg+3TeRYCrlPVl1IMYCUW4j06PzcmEhBJOetiUA
vhhLEbOXr1SbUlwbEQjxqH9o/KCk1JxHHuULQ7+3qgmkJ5ICF/iJrwmC2YXCbOCt243leQoPG9eo
x/f15tXL6PFlY3/jG4VzCQCFugcE4ldKbHF500uMXNIZxSEorIk2aNoG3VWJg9JIUrqIThq56nZP
sFTsADiDIY37rDi8Y1hSzUkBIhRAdupEZhV9WKcBD1DxtsEI5DVwfH309iBEgfebdzO4d4VGUbCm
OOOU2xUQvUZuBDLx7gIbzziKnn9eJFkrZyUBKYgF+syv00f5X0OqLeQ67a5ajrvesdLMswRasqwC
yPsYL+Uk7JThdZke5VIFLtewEuqQQugSFT8lCSDxrZijvn5yYQpeizeFUzb/YyiJJu85GNi23KFt
25EmbcoMyHe1IetcrWxWOJ5sfw3+YUsccrNiOJPeAUcUVqxkoZ19wD3SKwTfUjayNsPLZRntqCtw
rh674N3me7Ry6WJzjII54Qj+8HDUCxEySnQUyN9e/+uDLFbrPxPIG7VpuHx+AyS11sARKZDvvcgU
8BbFqiz9ZiyAQVFzi2flPt3P5C4As7tLlA9i9e2EVSr5tnBvqI3ZTNGee2V84Yevu2/0cQdMCNoB
iW0iBBBdfxJHhXBnEnjC8Ys9FF8pbGYxIQZ/H1F46ILj5fU/6gkAagBxwOn872MWz2iaQk8tXon1
BVSZoFUc2BK5GMAHcYOLdFl4XuZyqSR35cZ0z/gTX80L54EUnsdxhhX38ISTdTIOCd9v/qQDwsZY
rcIsmsqKtTZ4qOZ1i9jVrBRrwyEzzKmF/yIQRC6vqDQqg5LheA04REoVxaw5cgkZprHbOlkplBGO
7VS3qB3NwJo+LWaUdN8whY86yTCZx3DlLOJwSs+viC31EZy0gY4zN85GMrKknekjDb0LTTCHehfm
F2fBmercqDbGTZe/SswwMMNMiMyQF2wqOXnvS7sfU6OW8ISfpJnoUGKamrkFi6orjORI+6PRShRt
dL7zO2NAuz+51uaX+u1UEBzo6YJb0pMvWsQ/9NBYXnXPp8JOG7+A+k1aqWPhfJLrsMwAg47io+aC
rzXB62CrKCKcIeNhrHvUpU0wo0/mzfOS9vRM/hSi6LUWZKwadHGnWNUdMJUl/T9N/Xoxwbr/hTgf
ZamBirCZ8ii9eq18sUOlqFJJ8x98jJn9Zwtji08O9Lo2v/LP464qp7BBGnq2+Zpjk0XybcTeuGUB
74BdlIsJM2mTCs1IqexcbV5L0SKz/aky+HIOQBMWaDWmdP2sig/bHN/ja0tvOlpn77p7GUmuFsB5
h9TxzGelpM8ZSFrYZyJrhD95TVcuQZQzv1Mis4huU/azLJvLdGfpG2e4hBanZDXqrZO0Vp4QgkFf
WDWrOhBxTuBrVLcCB4hnT4pkcCg8vazLX8Hhe2aA5SwecWC1tCL/kowZpWdVpyZBflujeHwp3Tz7
/WuOlXmZTaTj+cvlHE3gE0FU+qbq8zbmuGOPeRxh2jX/NXO0ZRZf7Ch1RWXdbd+3XQ4n4048kOYN
aoasaa8e3Du5+Xjldx/Bou6Vgutt/QX2n/XjcLLKsGp6c5GuUvfLrur+h0OtvkvALkrPmdkCkj+9
cSY70aMmNp/mLMc1dJr01unecjEckGVIAW561GCmBuV4sdzTqBfqID+Z82UH/Pri6Y+z/gOgCu8p
y613DS7YEiJyFcQvqZF9XNGvTIJOBpgfFUQPDZ+CJBTIP2cA48fx7skL496tfm0D90uXCBWobzp7
3HEEuiy9o4k9TCKYc02OgtILnihXFvNyteCvhrj99LeiZEU2tN5ZLsUSV6hokfragyhkI2iBw+oF
GOnReZouQQtlQVVjrCo18w6QM7bZmY5/JGSGHNZkc5Ip8GZDCC6xbofcZ022ipsvqkLMq9/KlCLA
/o7BIOVCd/twpLVJA+jSperHNqp82yY33UwjWTKYaB/lqE1feRocx/7D6Uy9541sgJqpVFzrINzk
9ofBf4o+oeTAvMyNAlG+X8/InoJBYQdLsUgDUSpjQguEu9WrwljTMnbUIZvFSpPRxxwqjq3d3T8e
6vXabCpxLBWsGHlHsoWGu4Qps+HFQXl/FmZ1jOg22glQw7zeQNbG6xbg7LeEhEEmPVEEdE/oKnvf
gyukfAtYIIYsr3Hf9DUpsbzDOfI8wuk/sRMveBw6H1THnBqnZJnc+xKkszyx39/GHxIeihj80w8/
z4VrF+dgGTUoJtD36zUGmRGukqqBnswLv4/Xj+32V325DDxNY4N9zC3r7jlo7woXWWJfFUh3n/b0
Y7dGrImeqdbqQlaYqpNichTAeJgV4ISkPXrmSjmP/3qRUHIQJumvSgTrCnK8bHnXSmcTwDJXW/Ax
onAjUjAyezuIn5lWwGLBmEJGkzYI0mXo3FgUThj3g8BBWngEiHRfSaHst6VxqqtnMcjnCBJ+aqhq
NX6vLHbHltZwrCZfxS64Tc+Vd5X/gRO+iKK5752+TJDeKeVbAQ3GboIXrZv1hq0ORpFhS1UN4q6A
1LZ7aAYqUt7F+070fmzoUhX4YH/LH4in+w8VgykHBFKraf3nv8Bk4REQ9ryz49zJkkmklwdmUiQX
FLS96SOFj6B10rjhAL+MWACt9kalNYHR0JjsO3CBX7SrY86RBSCRLS3MmhbZLEn+Cbr1ks0cxN88
NQfb47hQvbOn9TOrNVhOwlG3aaZYDgY6P8hslV79nuYCWz+VBRQmW1PnQI6V63YDG93JqjiNmfAc
bppCTFm96PwtmfkDZuFzhttI2+AX7IG2KYKn19GXfvJ0FzIrBZMDzvxkdzhKJJThmTy1i3JBpvbh
2f4y4CraPOzz6EOeMzn3COcQGS2XSnqO6uDPlol1L2jAVdVidq6SWyJKPSeRFkLXBWzj7kvAquaF
62h/5J+zs8EsThD6crtZnEkKWKHeogfhOec4K+khEYLkW5tp/kKdXpvr0oPN+U+lO9v8MYfP/+UJ
hhhhLhW96QtKxeJDFR0MpF9OyD4tVzP1X6awI2O5V3zb/hCNHyXRq9GXsTqxSoXFajThRiHaGWY7
0Nn+Hydy06zcgpItsn77T9tGnfcsv/MGsI16GCi+wLNf0ybtDOgZ3gZZ078TqZ2SW52OFw5FCh8T
R72ATv5G8ttqhtehQAigpETjdg9uWCtYOkpMFBtHmqMJvZLgz+geoAzWtjMTIHjCYL1ZepHpn4+h
Qon1/pG1OdqY0FqUUn1i6lE+84l7wNAwDF3QeRI9MnNEMYqGaOpV5ej0VOTfeSq0MxZkJ9tsdT2K
RpI7JdSHNihiAr4NqoOOKERZxtVWDTbZZDmlleDBi/YJQY+L64LCv4rzPaASKaYUtAgtuJB5Tdh3
60dC2RQeKF0yhlrPjEQ4MDdLFKKkqgAyacKcr22R9YI+mrBWSHJWZsBZzJ4vYNSRDXpmU00EPA8A
zlrzMB3y+ZtCunpxUY+2oxUPehAkzSQ1YGZD5r3As5NNWpqfJ66+Ktgcc4JWC4N9hW7Y27yqRSal
kz1urCTyygpBX6e7qTr5WuXU1tO00QVmHnMHHhZR+JAsjOUKsMB1V7j/1Gd9DQVyWEPOCf7B6UyS
154gpXKE/v5ZI0oIlptKffDwmxCfjuFyLYwVU11ekNS0mufmb2zvg9VcGt2BwoqOmVXzPbUqH/lu
dREA0YoiuueLmg54Hj3JwRF2XoJKYDks9qNp6ezAGhgLis0DSO9hc1CSCtoaSMH1mO4csb2ggzTP
gTGppWZZb3FZWN5PylKiKlRC1u5lexkiQv2V5PHQmC/jhV+ioVoulBCkt6zWUYWa01DV3aatd6OZ
2xigYV5zRH4LluEbSeoUG9dwj2XoUjOMcGBAOmt2qJ4IDjx10lKkMw+NddZH6flRtececrqv79EW
B+5DzvsxVZweYG8mGdlpMMwJXXYFL/zskoHvvSOozvQ7lQXOAY9t47kC33U1pbZ7EopbbbfHceQq
F+XjOyCCB9uSe13hVG2LgCJvFI/p2yFi/QJS7kBlIuLa6lF19RF2pQ1Qb3GRSQyUCIsIEgH299+t
E8X8LtqyTM4PPmVFy2GJ1utiHS9sr5viRVFIPtl4FLds2pFhVZtsT5DVNlACkgyqoOtRxFrM/dH2
8GB/URWARsxVIAVJpveJMlCiJbIdgcgQ6xK9XNi+3f0LBwbrvygHJ5clAhnR9eSi/VSOpSm0meq6
QF2wn7CyJstpW/ANPVBaFiIMQTAAHEunyf+j17GQlFvDRYSJ3YwFIfqQuHkH+om2Dcf7qMGojt98
rQX0OqeQNgLbbn/hB8SuAbIAH2OGd1b2n9yHFNPbZBbku58tKd+qYJX9mm+fVVaoKWQlW6Gkq9Hb
v3q7cQVLriLxWOQYc9TNNKKRUipr2jkshZQLt4GJIHPdjFsgf0tcQtUuMwQ7FwUVKA0OZIHfxa/D
NfMbf/kMn4t+8nsyp+1BQJAoMhi4curr1clzk5mIxrtDvUCrvM4rnxmEnp3pW5ZigqDa87LcmAZF
UC0zjqPubNw+MTq8Gy/bzLIRc+8/Le4GJX0XfWHDk5Sz+Mh+xUdi9HSbub1tF3rKBIT82VkDo4eQ
ncb71U5ekJfYIqXg/ZiLeArVyUHBODAWt5aOpH1f8cUYPT/2m2bTHx4V/mt83SgW0goz1kXRvLs3
Nh7V6gb/hBG800zOPUoZ1t3gV5iFsCqeoRFtuqb4BlIZuHMv/PFzjeTw7QQPeg/3aR10bEtmchBg
QKWPw8PPnuWB6cBDjvZ1H2166lyV7DlPxg1+s+BHana9KGHaFeFmvF2RZA2LeaSDJ+yGWUWJqLdO
fB7Id7ToV51OJabTjfG/kMxLVDNRS2dPojrIO1iW0u2rSE0x/oeRRTXa+A6bchFITCyEFaZVopft
GU/EDfXUH7P5l07Vx509XeAl/dHx/f6ydYDjzUf9ZxIXKwF29yzr9wHZorcAvBoFA64Z6gwT9vx0
mnKr5GvvxfMz8A2p6Cdc/PWhWrPtvGzIOaribOfF2IQojDqrrMVQA5A7mlgVP1kP1Yex6cmWuehw
jnPY8llaSWLjnIG4lw83O1Na
`pragma protect end_protected
