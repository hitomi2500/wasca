// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:20 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lPKCd57RFUwqf25nFn45wRbhlTmTpjZX6gzNZaPx5xvRgMvZyahGyRKsB4olCgAX
l4litP9KyoZPjAN80UqjFQWo0qRDl0WN9RkiUsyof/QLYAgZLI5M7c10nOmM/oAx
GOfz8i0SmGa4tAXFdVmA1VewJABXjkkZ99FLct2QbLk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12448)
1aCf2eNyI1LIuJIMw3bLkOvUjN7lPKpW/0n/1jah+IU0rYDJFjP6zyGYEFy6cqS9
r6Lv6VOo/Bl9gg5u15DTxob2myYVBKFMNXFat724er/uX7Q8Qs0kxADug3V4qLRe
feQloymIlKh+2A7YLcGXT5UYYBnnr8498Z7dRwApF6njL2F97VnkZaEZ3KYIRRlO
Zms4xCg25zXj3kX00bk4S74+tR4iv+GuHDivQo+mc0N33QK9hb8L+/JKK2ZKPpiP
fe7JTwa6a74gtNZT5572sEDdEEpxqQJ+nhjFtPPROA3B4RUKU8xbYgP6IPq1+SDc
dzrAsA4yVeJGqV6rV71yyRa9Jj23F/azoOJsFhgcGl7jH6Lq/lzMDtaFIDIqnoyS
miRVLbAE0Of5eodjKWx4StNnU7bjnMhH3UggIcR4501Qw5G+PF4IFYlzJivE4omr
/oMIpxmlS++mQGfl3RBb5ScUCzCJJ7NZ+3Yke7VUtThp9CVkI9LL/b/u3Yot/ZSx
WfjOtsjwqGErkR2nHB8LHv+hfKrnSUvgrOPb01ez+lGqAaqifwMDKVPmxpYw3Gx9
1Rqwmz0iyj6FR0sgnSRs1zbl/1F3ifk1ByLga6JI7SEpUS9Z9GC3ly29oLrRwo73
PeIMstVEFZwiiGDVPi8/QCUNJl3jKd+skZBFjW+kPbym0E1rbVfjptnT0HCZ1Ps8
p3uHPm9hwGxNhTrOBLCJaoxk0PIVyebYWmHb2MgnkhhCJOgqn1KcUM2KUKN6vA7x
tYjyh5Ed5EdmlYNqU5VInvLo5h78shymo/Yhl9JsrsE5R4LsGBrGfalUQG07Bl6C
FFBkwfDRzpd1KIPs/XsfLKa0xRCWau3U6us1as8s3dp47xdPsu9u5kfe7wNRcdPn
7lwaV/ymwM2XAkXK0z7mLCyX4Lo5pYrUd77kQVgGXuJ3v5vSfx9I7B/iZLWykyw+
jpeCF8KjGBQ7jpkVUR58yfnxBR2PqC5CgBDDdKHTwjgeM3lXbiYPG7SKs3ish9Qi
61ttIDYOf77BJzh+oU4KuAJaaDYcn9tP6hU/zSreA4Hz4S/wNoFmatzS2/wKSJV1
SwuPBI2g2ABriZWBofUBUe92NWdPqaDmUxnCQ4940fSWJu8cae5B2o+gAwBDQ1xq
5dlm0vvTxiwqw3GVU1/juM7CZN+pXj2SbzJBBTFTIj37lDnne/70PUy3mNUlhN4b
ik8cOMysab8PjAiMOXftxIeXZC0LLt3BzNJ64CZo9R4NMqJv/uYPX+ohYbtdpYCl
xmASHLqUwpgiOYMp7/v2v4FgCdAGBTRCIq7vaH5aVTmtZWjEmGs1vMIq6c8TM+nJ
2OyF1VZF94jzSOnBbvlEHLrFDWxoFDJ5unJQaCLvCgYVhl9PwHraLU2iX4WTdnBK
32K6fMzPpZ6j0wPlvplGtG9dCKh+eiw0aUcFUspxSfd1PoHGwcZzX8rlGO8+Lm8d
jc4U+PmNt0NZebZtpP20uZIfN2yy4yugjX9y1Xo5hZNl1nWEbty4xFJD5e1+lvHk
unM5mn0K0C59ywPnMg8qu2LkJZe2K/+2peIZ+gzOLR3Fku6xX2pqzWlIJN85sOD+
8M+mvogSuujmSSr9F8NNBkctqdyHhRH7BxzFGxEizPhhFoTQfmuhf1s2H8ONjK1S
T2fcSj3ufZXSh0J1c+5pjdkW8SZ6JEGh215NI9ynU0Y1kk6fn9i5ZaBT1m2h4cLR
K2SVbK8sX6hBn9dhxXY0IS5St7fZBZIL0654JKbrHjMeZz+uhysbDLFstYN4OzOi
qifWHTt6JRpnPOYqBh+I50OnYD5V0Iuv2HGdq3IQ3IzhxKRoOlWve1IrE4V1/K0+
3wm7jrM5EeHe8g5LVERaYbMJ+O6OtJf3CwWUKUDIbfEZtJ72NMeW24Flw7TGzxJU
DjmwoHfjRGVAx4QkDPrDKu+U/7+AsjtupORsGshBbnmrs8FN/fBZtN4Yhf79Ty8f
KI9qpMlMgdmJstQbp/Pz8CbSY3Ksa4YpXvtfvkJbhc1RUaQCiAZ8Ke3YRkd8EUPa
Al07VhmgJFZdBIx3KMki2gq5u/2zgHhu+tqtnmwjvhHIDujDeyOGKJlgBBRMqg/S
qyd7xAofjfXWiMxd/rKH+GgqGblFkLeuVjJoADjNSr+ge6Lu+IfUshjy788WwCpZ
evaq6ZPIE0RFVldmMKS2y3l5yhb+cpoPYGvzFCuY3SMUFIG2Y8NNeBtzDPiRxxpA
4mlQ7wZsoLgoprEre/9gPjRg735h6qBVjjmJTwsfz0BVGRkxOPk3VYPT8eecW17x
x8d/W7krRpILrrAW1BJFtFAqyupM0NbJ40c68LRiTe/N0CP00tIo8rWsbCqjAzOC
C0UdvOJtCc+8nhmk+GMyhAzhutOOVYMZwjg08+4y7FoQhhXcKuPRtZ9HYqqN7/ux
vLlck6V30Yuj0MzGmY2G50i07gOAZw7fjAmujgSd3gNypNXrZhYdG3sQMAqCUmoB
dyolBPVBtKBs/NeMwI3nnWF3llH9cpcos2+ASgvqBY+YZkPDliX53wLaMGDd/XbB
DfzKmhTYvBuXQvFNBNQ22q61ASM3F0G1c2gnHfYWd2k+foUlCGyYCKdzAUFgt1Jx
IP2Laolrhg0+UWbjPZ3/dWv3BNKq2FwW+ZIPL+hCHom4uTqU+96cQqvaMAZh7BRh
dUiroN7rHaYoSPBaw09ppC0RCm/eigRQjK45+dio97A4HKQH+xxvvFFWMjS0YK5Y
AAY56VV7+nS1QdjJFQZMfXkZq83BVdLTg5LgSdLoTm0ImrT4EY2vGpGi5jOJvZ68
u9kRtOoYg+s6oinCUD65Og71yrE/G/mYu1efMzecWTFbm8lHVY/CSBJQnNGOCCzl
SqBXJXOyHzr7umaDqkZAHaYyE/PFSVinlzkl9YpcQLmz64CCzHAG2IxoWlXwqMlt
QTecAgehRjxxYI0jL+RHmeVGvwJun5fc/opdqqyLKglMSPe00Hr6ypLBRV0bgrmM
7/HlB+s8byQ2CNQMVkWq1gnxc44F2gOet49ugmUbmVViiY41q4leoY+2cl/YG1tk
11DoKKUdrxaUjGKRN5nrfUwl5+p8MytwIAn/z8O9ZKql5USQRdgSFEH26LVlbgm9
l7hzn8L4iwn+KV3tHgRFemb2jakFRUgY/ho7OqU8dFgkOukbYpvXCMRjnKiRuk9/
+PJyTENTVwVOJajHmccXfb6WF8VMSyK8GlweIr6IZnwXgqSP3bDKSd7I5mOnF4o2
JVPzs1wY8+apC3fYs4iYX701IF1QgWo+FiZQpCmgKPkXUuwFlry1p08Oad7qrcFq
8C3X9oi8r9SREFNdcmNgy91vZUnBt/fNem2RQvOshE0Yrx0DSFG/DUS4+w4RblcO
/sL5T0WlJgT2T1V66yuoRjDEzsWy7UxBzHe7t4SpyHOaGGCf8YDB/oBDwZCe1WP4
b6C3DTMGfjZC76sxA0S6NO12cdr1dCWCytr0XoinAfTsG0JwDMXrnlvFNSRt3G8J
5g4+M6i73cWbeua8T8lKLtgC0oquJwOqRKvQVc9xksiJqOIQgzLjnrdTjwuji4VG
w0YFAl+HP+g//mml7x8xt32kG91pXULf1q51XmHD2cEOfBSiyTS16SDzwg0YYjFP
b1a2cJuGQh7N3XzfxEALw1NSNs/LhAzApOcU5GDVwVN92gdUd9NCuNoEjmJqHslY
sdT/dPqk1RsX3hLKInF/YrBrZBdB5jTmk2hfD1jgQ/Qqzuv09Zad1PYIouaVMZSE
NdvzTyJ9f0UBGxZcPZJ6DTR/roERhy/IOq8KcCd6aGx+or8GGa4lf1LSx4mmiwg6
rNOdyIoKPUagYggz77Y0JT5F4EpfN8wzpZ9sydlTBgb1iTtqypedes5hlwUvi0yE
HKqq9qbkyGahvKfsg9bAzO/Yz10BLwVROuYz/D72WuP7DdvXiB/aC1GpU0Pl6ZjN
zm0sJtCRVUERRYcWjxFVLkFiID7Mwx1oCrUA/ofXoT2cpU2P1L/m+eMvjE73zVtB
PdNHwIzYyx2OiSk7EB7WK+bNKmbHGDjZ9az8VfQ5Cle0InwhBBlJCfE3s1LU789/
yboahNAsCOkeADJRn3XQpkRdoUjIxnGQRu19SlwLRY5Ii4mO8/8SHvKOHa4FH60T
JQAxUXTjTdoPyFjCzyQVoVgE6l0SAartXal8wv4o2/NQu8dZEYfeunC3cV6+DjnI
tVz+YutFfz+0Cn4Va8EzOEuFFNHcZvVtFNiI4TsT2s3vc3FF3k8pcuc+vhDJYm0T
6PShAd9BCed9WLomk1NQNBCiExikoNwXeALZ3S3RNJgdAZx7BYTyYjvn122tDgLy
RO/OJUKpPFbub40tCvyNRITcColIw+e0WY6zUNo77HboeigBGTaan9mchy1I9YF/
16A6Z6H5a0/yOrAXupqqG2Tt8a1KgTrv1rT4JIUcKYDTqqrF0KHpRBxGZ2cIRGxy
5xiU+pbj5vdYDSt1emjMExVegQZPGDEeRnnFLm61viBN2GUyhbU5HtnQ1a5adbmn
IrO/DkyNhT5FCemX195YnJT8vZi3BOMe9b7pNIPbhXBrIl0p5eOPOnsyv8Zpss/r
jhx9pvMd2nEJiIFQsUCWvSHFbO70iq2c/gorSOhFNA3Mn8jN9ZEGjj2ZWLujAUIP
8yuPobYQXl+IztfgBnt+dpQTgcqi95or8RllMclApsBVRcfLbjlaB3mKoHfvAu+K
fmXM+5RUdceTp3o7lNmi2EgFJYkmW3sK/0uYcEB1lhG5fFdeJON7nTMHvaR1Jk0W
1XwVKRu/gEp90zTpefmIGDbLGHRv2IWSKZuevBDDpWJvtO/dx5O9QKn9kvE8Rgaf
t0ZDKT8CocM2GtqbHLZx6Ai/Q46IYuE7/vcD0D+RCRo0sqR/dKTEhoelBK14XQPP
mV7Hneni93yTMdOtz2T331p/MkT9pcjQKq4vNpYt3p+rRzsiF+uSWgYaGZ0fC3mn
Qk1+3FMJZ4KmoAbvED3XaXIVI0JORNVWcd+8GTcWiXeV7d35KiiOOhxbRR1ZTT76
xe8R1CywIAllLH75H8/c9eYJLk1XjHggJu6J5hbSxCssmUBCCykvl+JFjzZR6z1A
YFkM4Tg+XIoFS2lG+aIbT55Eq7tFVh+9aBXjz2VgSXnaITUwOASeGmpmE4S0bUin
ptj1YGeF728gTKAKrLSMi9KGzdpZbda80Gce4w46QfyC2zjAbkv7riymJDsAX2Vk
zme2gGnvYbUOToCnC0Tmv3RooTDzIWuv0wzzPl0rXfvaoiaiZvlQIRZVsQnt3Kbz
f75BZZ4gRyBljM5FFe0BmbtAyTXX0ythsC9ghIgjvODlsF2KsaCXrtlzpr1e+g8q
SEfF4jhmcMXC8SdOf8o/kPz+2CXYaVe0wFqKJuFvrMkVDPav9roLY6aNnMTAKL0s
UrbYw7hya64Lb/WkZZiFXv5+61/ULIRvXBffgJEPN20qcfwicfvIFa96kFroJ14D
48mn1KXeYBVBlY05ENtWWYcxAQaP5+FraZQPzMIDzDSxknQALpYwfWq0WvfPPGJW
fqWj3cTcS2dC/oBIXETsPeHDF6g/HJT+2FAUFRqBqgXePgwk8RtXL6AYwQlzZq5h
/OYocLl2UaEcO/erY6EEOgyPy07Vwg5zRJaX3PsXfQsN8YApvu1sPOWkQr3aIgGH
ES1K7Rksnmn3Dl+pkBs5RNFhMem0e/lUB0THRJ4H8Utg+vmK/QGI75JKNt7DUR/7
n523Ks1HCvg8UzVDUNiigVh02oPt0c1TQ3WXiAP3iJ2LcNtqbTVMGWdNglnLhthq
EgMT2o04OwZXRTWidop+8I33Qx5/ItlFCD3/CzbHjv2sYN4LCXu6HKoTDqgvULOk
qH9uZjxkEEM1W0jnf98Amfz19FeqDFEoylSjYKAmBzAAYLycVsOaPVrbE5D1g5Gx
6EzGSf9TDTiJ4uNPVF7VbR5FEF8oOgTi8Yk4NJP681hjSpAkmgoOKK4tnVy2JhVg
sC+I4D2RPaAiR6DBPMPfglD8RXDUIEkCeYkpdU6t+d6Yr2lDNDkC5isnqgxAjy7t
Yn6JG6CrtfDvVOTT64TDzE2wDPN/qdSRN6hknsfuFGEgj4PQnekGcJgs7nnF6qAW
LLe4LjBriyUYPlSU8Q+E6t8LH9sGL0Y/WMFyNJ09pizEmpQV9YqxRIjxxbDIeixp
2edvRq2RRLTpt30eWaZ7Pon0TIJa7j2hhTXExrMesyqQ2/HD8tZWlQh0AWC+UnZ9
iy9FsQaGYmYKgM00+1H71C6A6hOtdgcWIHwUTpRMLj8Q2L9z25/NEu1+mrk6xzS9
r9H4K7He+ST2MwYrwWvjjJexS5bzYICpiXPHPTKEyk4O16Dzi5BJGlVJBWMHqggb
tj9p72nVcwvGLohR8aMM8LMGicDgdsNxNKLxy1wZTNKzOv6dQcjnw0lCsxb/i7KU
p7Zl5u9W8dgFQjgLQUAE5vMDq/BRhc81o5445QeNBdu+plX2V/9ZslVwB1mkad7G
Q14J/IToDqpKO3xRI3RN2Phf7CQl8u1ZENs0wAtlvyDDj0LMhqPC6I7T5DuwTfPY
2EAgK2y0/Oh/dixNklh+wcy5mfKJDUbcKuftvWfhsFGaABFqyTN5vgD9XA3cQrwq
Z+iVZYNXEROrEuQMKt9/k1vyXwpeZNUEk1jaWzYo6G+MG0q/hn79KghVopNV1WyR
FZCgOXd0NyzUiKUt9lH5cAebbSP0rjdllYo3xPZkBY3VIP4DlioqqzdfvYH+cUda
ZSOQm+CW1P3j8Wu2PQeciaKJP0LiSiyJ7fQsuqOtDjzEKXT6TvE8ZqWCChW6jlq+
C3pKaHKr/SdY6PdDX46f54DDZ0xUC9joOjqeVMmfSqwjINIZhmomomEC8xY9UPZD
LXGRqozH+nah90KPeFmFMhm7mkQ3XhVccCYMRXRTnfijccNUraW4ir86HNpnCsiS
QEu7nv1uVo2aPPLklwzBAbMqryySeXptV6/sDgD1sTDY4CAx2rQxOE+Pjf+Qmf3F
dB97csFJQG+NMB1lxCduRXW/BravZCiP6xUFTyU6ptnL2jEz5ttiuQP6IMLlG909
2B88n6Na7qq5+75O3JuA4w9Bn5GzdTnDZ8K0herLVRTMWHbOOJsLxtHn0UYXXdEv
24m7nZXmuje2CAuAD0xqa9zKiwuItD2wFHLPnydqIgUUvwoqkFbZGyHxra1UJL7B
mrCs3pRLEVZ/k7R1d6H29xj/BcGWOq9Y3u5Duki/D9aIxD/3Qn+nbfrzfMybBiCj
3e+6d0EmlNnBLOye+FkORYThfQTX+q83ySZtj61d9yKSo78uEpvj0pckIVSVr6B+
BTwDL4+TVn+dsyXVekJOGMAgksOOOtSwpWCLGsFQj3rLjmBlxY0uqvf0Nk8OqnD0
9wWZyxZI7W4AmaLTDc13gE1ktmqBrdev/Lf6h4W/UyzeXAGoJ7oFmHgqiGkBTa/c
JojeyWMpStCLgu4TBkOTAXBthp0lNF+yHv4PT4EuYQz/1Xpurd1fmxMb5PR5M6ep
v8eXa/cHPcCVfB2EsQguV6tfKj3iUWriGtgMrJPrH2KADxb8SRlOPG3PnbVqbpJF
JxPsYDBgdKzHntgHQ2NvRA+xGrQOZz9/VNlWSAK+RRjF8KKD0up+/tpuf+7ZJi/Z
1oooYNQ3LwjNvPCoGikgOxg8J1IiZGP0aDYzCn5DZwLBU1NhjnrIXbkBttD52PCI
H0h7J87XlkNQYmgOnstKpppv98qY0YUZF0xBpFYcnPG1Z9FsAlFZ2EB5EX69Ubh9
czLudxhAD6aEDxWa3L7L9wsinRAvq3V3xpGDqxkOgI8s30hfK6Z/Z6s/u0pPotuA
b0QGOvJ9YXRwlNvJVHhLJTiI8G7gspREb8fRXQo1PFeh8XdjUPC3eZFHA9fqz/0W
0pHOKWXgtELVCdZPbz9rsmndL3HamOrYngZxy1RCe7ec9ZxFchrXssB1YqZoR0uV
Rb6dZc8VyBw81yO7XgncKZLw80ytxWQmnFak6kZ0lw6NS+5CTvW+gx9HhPInSU9U
loauN4LlYXY8JiFDlQe85w8AhRna3Lq5HJdGbOk0IOtpPsN5+28yYsIP/+EmjQz3
GinAoaCeHDAsv9BWqYQ/QpyAZOAVi60ZalJEI65QRbo9YsN/lm47RnTjn0oIJDZp
xHK4YvSwr0Siv8sGvI/HAs/r+iGathn/np4C66DacNxg/GSqPqlr3wV9hVMy80Qb
rGiIr5EOqzjY2tn1M6G6X2MwOVWvYZLoEyqIXfQ9BC6AO3WGMqJOFhqB7KYlxw0i
SmWib5PhCkAQD/K3DbYkcmfvxmXZ3zLejQIfmUoggyjHDuh57kMn+5Z0EJ3fNxNv
zIKO5C9wM5inVY3oMqn6vLUOUOV3Fiudq9IBb3sFnyp9Tgdj8IL1EwfOs8ITlF1R
Y9DBPbkqKIfoFWZVvNMf5lQY5Zn7b2b8Fc4BikOxEVJcUZ0FYHFxq7Er9sY7rBhM
fiFFb9PUYuMAtNeXwyqd/uhK+TXsauVDHIjdaCScLrKRUGzZAGX/z3Q28JUsn5ER
3alw+SjO/ZHcSwB41GPs3h0mq9TH0AbDdlknkmsAieP0/hAk3nUH1IJetqKcCVRB
G+yH4Fn29ymIQAzdEbD++twCfSiA6oC95I181qlpAY2zQrLbgAMy/uw4D+f1Ub2N
XWMu00UqUhrmoaexYOj58ooHbiFtzmNkEp4ccepjw+30csFS0WuZG2pwjmCiUy91
MW5nv4ICCWnAZKoOKDreT1Le2+Cof96M2j7piPUfrkV2/5hwoxNpG4a+NGIGU6UP
PiXw8VLGv924zVxFStbJghqKMkcpxikDuKEoy9BQTmyiXtU5Q/EC91FGhhIzDDFw
GY79DcwwyG1JG53ocZiN1xos2cSvQmKzYRWKZ7GSkMoG705Xw/LyjK5T37l9BBOg
h1E1EkL7WpBDdebO1PlS/WDQGTL0W2F3dCQlxlzxsJ0Qo/oaOMo3390SwxxxB8iS
Dvym/DLLJl5qP5zfh4HatNOxCp/r0zjH0M1tPtOee5j2iFrhs4f53a4KRCq29bNh
/+N2gR+CXNxVLTOsrI//p5yoQsXjeN6mEjnwg/UWI4/o9qJtS72qfWcmbnXaW7Mb
lbJy0ZFEmQ8hwSapJFR8jCt4sZFqy71zsylIM8IQR2uCzM0xjsgPpZKmUCTJZqg2
RQR64QocxpN8fvWI/vWdXgDH6Xs4vqs2NCuFGVDjh/Sjr90GLtiVVj3Hpgh5Xfhz
44DI0kQK32rVnZTUccWA8BoCIObkrbnemHnblVp8C4vKJVKeJw7VbATgk74DwYXN
pK52RBAg5dbADjA/efgN1OtcGrjlZ4w4vzvab1eeD4ofMSTEgivp0Qo07wORY+k/
RkJUgyvzzj3+GR1ScKLnQcKXvnpY9ny2JRIkH7E53ZmbGuZ68sxArdkzWb0r13ho
pMOxy73BB/Qmq9OI/KM7pr9RYk0kFfgzQoVOHzBOcfHiHudGEzK1hwvuFX109SpD
PFS2p2blEaVOplAAeso/uC0YaKtcmC5yACbTqzbgPyRwxcMli6wc4VA/Fz4ft6EW
Z0LsWG8yd4cLRLgeShSJrBKh8va+5/EzL/YuLGYO55EVTwesapvUNarMXfLknbwq
+pdgMY9zSI3O8rSucPIdJki+wBOktoIhUBu/UySyRU52QLwyRT8SRLIZrdNUEyK0
NhyhtXGZbfSX/Sm/p41PxncnK/b0GeB9rWNCeHB5dr0vZy7kceQFAAGSXjO4oCp3
fpnYMKvuy2jpmtG5+OhuZtABugbE7BLQz2I/6hWCUCKz0OtbDBgMbDoXoo8nx6Md
tlmZ6YsFkbrMLZ6nqB71w1ILDoopVcrqRRtrNsG3V5e7v/+6OgroC+QkfKFGnXJH
vxZsviFhADDv/oTfVoePqmycqYxqsmafYc9EgXpO8ab3DxS0+LRmrBRyNPX9JkOw
xF4VmsUgipAN9O0UOItr//tdlRpen4GzM8ADFSeZhQBj2+rG+yIRiOzRzT9osuO4
lj90tVj9Wd3ETu5HcBN3J2Xj0eFo1HB6O0yD2/nTbY/+brId+rTrLXyk2oODJOTM
XZgHIDuFQWu/cNZe8mftZvfQDDXn4zVv+k+RlgPSafOxnDCMBtp8ZdGjG/LFLzNl
VJWWyjPbNcO8JUXb8Nkg6pXqX8ImgHJlRnr1svLbek8gOue2IbSkQmwBA48PB/ex
rWNvfyUySoXI48rFSzXHd2DqQTnzKXk5TpZEsunz/GA5oklglz2P9OCKaNybkZY1
lLrnVTldn8ueUl6mVzX3nrHG5L++MSsLAG4+C5nrZ5Y7l/e32hZCZ04RSvXJQmVN
a9KAvxa6qV1f4UH3nuJD+ubhTMI7uuQPz0HB+B/dkqazMykBxFGfPllifteBRiiF
z07j20isK3ne9qC079poivb2Of/l4XtdbwvNBejGe44VxUWf/uQlo4nlw8fucTpa
8YC+wuPdnkWez9UcPxgBVt2oJin9SXl0XcAwKxYd3r7DDBzoqUPU+Z9wOpjIKSKj
tnA3TFvGVYEgGdibatShi2vYNjoDrTFxqQYWxeR21PxRuN7x4i9YgeVsx4piASAq
3cdaualw0gAbqamAW0H5pmUVZRqma1QgOsPXrpl22ekexJe+xDu52KR7atOy1X8R
5WsI31Y32zHbjj0T8eaDCO/bX9/z0CoyuVeBxP3zGEBxLm1RK7MN9HnDBqcAAVFR
YW+FJxRGb7N9u77AgAlJYiFsapC+r9s/ArUCrhDLhVAEJfYA73y4VQaTHHnmG1ud
+L3UBrrCqEZC7o9wQu/Uc99i0rue0LElFIv+bUkNjwwjlNsdfZnhFOdtVvKTgKDw
mhXTGLNG+NS9aEBvOX9q7gFJdZw0adzK2ZVvD8+6UMDVmfd0oJwUc0EGkQB2VfVc
TSYeTKKducoWlgcvvgF6ZjA0ovKu0BrBz5lkBI3pec670tsbWWWt4hwACO60QXXP
ek1l+sMQCmuvyz0ty7SnQm+mna2lJ1BxejUOFh2UqdTe9UxKmtttgvyql7J6Zmoq
hhv1gnVdm8I3TeTGNlwdZnGSIpdh3TjY1WiVpE6iE4V7viXJe4JzBYkNdYDcxCZ8
zBZS4xyaR6xllsBSluM8J9gl6RX+32Wk+05XLPRNJHPetvs0C7182MDFlUPrH5a+
m9cmhsbPm6yJh4O/60tt/mU+uFG/uIpIOA9Xb/YMawAnV6FC6jWEoJLYp6FQ7srv
7KV2rnBYVAJxNy1RS8vsUlgsUBiStcewkcWU9afppP7op7xioSl8r0Q70Ng+GsKQ
JB2TaHIZkiLsTg6LSKndlEQv0/y6HaXIU9WjaW+Na+kSOCCRVsDzYjaSQw7MO2MR
xL2hSJVwMBAOTnXneqBeEMAplvA/s438ACHwFw9xtvzvnMHY99I3bF7v1Cj/VQTJ
uZ5/VwF48Qa7rFyDyPSjcRlIvuzRgYD3Fb67vq+l6MbhfTNpGTGEGAwwL0/GTfg/
rVJWQVPBuyJUKhPJbgRt5J++JPXnZIC97MkH7ewtaZC36SBE6Od2F8Bmlz4Os5aw
lWa4OjS8SMHfWKhQ2uWSBmeo45Wj1TotxK78ReCwWQEOMCL5ASm9q53nORSQ1y4I
m2hpU74rGGVIiph9QaCC0M6CnYGGvQaXYw0KwGi9OIDtQ6qT6RqN/QZ2tsdBRq2U
RNUgXCxFpLDMI0xtvvzxjKcy4Bf3YhgCXn0EIZLJh/z0q62F1Uv+/3zJyi6JlAn7
0AoV3Hf2n3NU18cDw1FvztKbcPtqN9v27c2e0p7FL+dTtqmegWJv3EOMjr8S7EbG
ElsrGF2NQwaQaQ+utLpVZzlMKnKXxp23iqLZX52q3OCHt6iCKfc1FtvBE/Fkifkc
baz8z8iOF7uq+U9QZEfBNu86Z9QJ+2beV1rRcr/4xdu7u91AyQJj/bR3vXQRR51y
N0ToIWlwLD6OIozZSWvkdMGFNFFJOiSiSOUz+0cZwwkZhMcBuTt8RSORs65+LtOY
tozXBrGQ7tRoU90BS2/LLmQx9F7pCEfD2UvsLZ/hFTeg2J+D3rzNeCflGFsw1AOp
W3p1OW6ZORc17vNhEmH0zilX2rqXQNSEHd0z2PamGSA01iBwF7OGXpLt5S03J4kE
xGlaTybYozWFu0dBYK/d8/jEjoIMgqYmJ2KNni5+HFK9cyU0qMxNQblzNreR5z7t
8eyVf6MFctYiyDAuDLKNBbYK2fO2Fc3p5FSsZCBjJpzBpVgl0eiO5smrDFsR4Hbw
Do6IgdfCbKXbRsBjZ7DHn066o7pwWo+BA+nIOse6FyAmt+gcD+r3OciwXrwfLA/T
p/UyLfI4U0mrN0hjBYRmKVkHTzfo4OEdWqVTGXXuUxvDTjmbZW4cQLoBuKOxZo/w
z7U1xVddtZzEcV0+pBgn2ljdeQp26vq5AYEugHPlwXdMiG3i0l6wPxZIZFZ+AWmu
WIuA563GFoSs0NWa3nhbzTysHrvSZsw5pMAJMYhu0ZmbbAdaTAphc/AA2gws2hnr
H/dyE57RuAqzmNxDie71K5v5FUnPaSb/d/+RZb/kWIn7IIIt/qQ71csl8dP0mGsy
7qrYXRTRlCl0/d3R29AxXxiej6+hZBDvzvZh9KOVWEEux2o7QoJhY2jRIpxiU/47
HKn7QqH30s04T55csGIqP6+MRwS3upokANuOpkLoFdBBu9LKq8HR6kxz1uEAInEa
qxn/NXgAA9IgN9ZwN0+MXW/jtTQSVuB83h48OImdBEe0tqYRskpsK1MKXRAvOcyL
YM2rpMo4Xfr+JZfwoHnOzHziS91sKRc6C7BS2ybc+IghmtxyBr17dTbyNapZjg06
PNURseNKd+FspSzDALtDrdCVF7g+X/baQNOlfS5QRkfUdBKz266JCI11twmbfCyf
uT3qaE0bTZlOevuYEWfbxYq0kHpvLFS4OD/BdjASTUBczQ8sQelG63tzKET8R1Zs
iRDtYA+yLo7WCmzeWavrvsx96VpRsMaQ3x4oIH3fR0WrxoHGaa4E4ePxyhYReAxW
HK34bTcsSci4SZKdOeNcC37lZ/Hs1EK5e3lqJu5pGGMbq1iC+1jbK7ikUR+eTv+L
voFaQS9jGSxv1/FUNUN6iM/l3HbuL/Z5/ydDY3ReWKKdtTv1rvslnhtpKohBeiGe
drlgkACvXKoYlcstTZQyDGBZtPYbEpNgJhNPmugNHkSIzznSwxYgJNFAZQK6Yh3j
F2jnHAIAPmzGlwWau+msc0gpPrzaJ7KrT4p7bvj7FtoMeD2zslG/czDj6lj/uEKd
6fNrTSZ3FGeN52ghNTNyzC0qLj80rPtnaAe+tXgsvsBZr1zrf8SY8lplATNrzVRS
/d/zLlHpwnBe2MJemEPyV4m7/PZd9f7WSiRXdsGjixCAloOUnT16IROizHaVss19
TGT8Yn8UcSJwbxj+eXiY3CWIZDn0Kga0ANApGg/rjV7WUh7Fs7s/iaUFmCGwml8n
macrmQ9t+xwaKtjr3vFuPPSaR9eXkme5WNxsqU0R9Pu7wOXe+/c/nYcdpvw1tENl
vRecox0AqXoWSBIMs4OQ6AiuuaeEE03RkuUSiImogzxbHVSEuME0giXZrs+lndyI
dqk4ldb8KrDfgdfGZNaeTiPjWdtfApg5tvqwLJmRZlC6BG5YdZVg1Z5QnLkB5+3G
h3P9IFFxSyBmwxNpQaJOoJIJGL4wldJ9S5lBT5F0DokQevy/mF+YGtThSJtliTMm
0qMUzqh0i/yj6+3MnItAthCls1OWletCG/L8PKHvS9BrJrlz30pUWvjjEQP5g2vx
7kXBnbANwpIdFJpbwByhpGkX2SSUozJmmu3Mu4CIbGiWFD2DEb5DzzRSJH4lXnw2
jBfPzCsKVFDzkXGojr3V9CkmA11RbLRib+FxcZoy8kCJjt4zvdIYa9mZLsT3XyNd
g335VMjhSjpQSYIDmzSCoDz6Wtf1SjJ4XusqTFZcVlZtBJxXSMkwd/MhT8QYGZRq
utgN5fO3SgDm8C9SPYpNPfYYk7blkdRerws1IuutD5AEtBIFq+++1DcWR1/TYs1m
8/n26bcFY6ZmBhyW5yj3X/D7GnQmhGBZh5TalKhxv6BTXdAihn3TTxviTaW/xNNG
/qOKrrsrI12PIB2fl9a9pMDUSWwn/mqaflFqqMz6j6LtxkX1ePUCJvwgJvhAVzWF
hqiNXMQIQmmYjg+k29nocPkSUfqJu+J4ybIOAgVZGBP6BdoCIebXo7yJ1c27oy7p
+0Rx6NmAbM8eZowbo1ri1J7NSjjf8vfisZ8aaxeAYhWNBQpHOmEuQtj63Z+9JSY2
Vn/B3NoNNBq6p6yGyX9FOicO+AxVviOVM5OwE+B4p7eyuCNjF36qfARzHf25abT6
HjOMv8jArkmq0Wdz1b9Zzpsqo/tIgfjKSIBgAIfWZcoZJTTguNvwx2QZNt7t5PdC
H7ltttsBcTkaDknryk5BqrXcV4eVgwbHT5N73250uq90uL28z7J/5pI219nZtRaM
sLQj/hh3ObQW7jJ8qkw6F6Evyop/p6f1ih64oAbIGm4OhCxf0zgMhcyzU7P6ar5s
NBnaMUH+T54Kuddz2tWDuvRPa7WypwkGxr1GExgonLoEF5kFvWGmCwV/bPEgCdbv
vaPnB/8+T5smpQGU49ePVHV+KpGYHV5RaTBziK0LdG5jjLvXM/Ip94COJY9DuL3H
yMgt77MNWDkJ5bwMeelzant2S/2v4XNYfubKkrZJlGG4wC+j4+vWjDMJoC82KKVA
cmLdNht6mslWUNne9ZywGlapigsbUNbNuirVNCWPNF0+BXVoMge+W/slXPUmb8DI
4SEbRXrzyduZ3traPtlJxN9pT5yo7302yLRcYdWKj0dlKPcKegJ+YjmRp/Hs1g7X
YoeYhKFX3LlBvJUtYVR9dKaRxWDRr0/yWh6lmJz5ZOEYf0KmvjEBA+0yIdCqb7pJ
WMdRMFfP2dXa8J1JoGa1q6Pto/T7ccMW6gmt+DBa+ArTQJCmke7VebsyPsp5DEC3
iLV7zq9vyJwiPwi/XGG2qW0G7YsIWHziou9vI/zS0MzTI9pj4/N3cd3yUnQu7e9R
nzQ4ui2YKyb3eb2XSRypcU5TYIio69+aaQPWCeRxDIs916E8I7EpT4PM6tofBccv
/LZv2jJQxUdb1D9Y3oxUFebkdWDUMdib+tCcuE/T+GK0PSgeblpQSmEUsmSYbw0T
ZgCllxYWqRQ0lgs0fXkeBThlsiCVv6SSpb5YpPq9ctK7jNwCgHQXsmrlwB5t4oKe
zwV7HsD/vU/YgExGfeehG8SPDBl3OKVqn81TbOplYOB16BPE4lxLpGVb00r8ZvAo
SgrgjJv1TLCT2Cqr44oqJITUMCr2ZL8qUehPvF6uEwngiptnmc3WucSxtkgSCMIV
JsL8NP7sST3SQmChZHcJ/481/CObqi+OpSqYKRMaBx66sM+po3ODyWMlD7DmO2Yg
Ie9rzMgURm/2PYTZwPVJJPEPMF090VMHTDkCa4/cumozp9WhbBV2MU4zjEyfc5Gn
uair5gAxGn5ZHOjAh71LGJbmYqufcA7krz0GGE050vf3Kb7Xd78qTrUa9j8bvpzZ
yd4fTyrd0oo2rJpy9wp0PCDi/OkN9Ve3WExNzLHbf2U7Chz/I6lUb0OhMj/HrMHG
Yq+WmwpcZOdS8gK6XVvKUSJ+omhz8IBwk1xO1aO23DicR4RVDqN5OcAIWYmFzVnH
rbNQDsiAZe8yg84fChMabEIufgGRkMpL2uwmx4H19UVoPPjH4CXezKIorKLGGSTj
p2qZmU7fHcwQ51Cb5vSGLJXonTDMnS+l1yBJpW3rzN0wHJVr52i8Sdcb6i9nrrbr
aQ+Ib7NyM0/5eOCM/TubcMT1ftLLTX93MKudV/6wAVuiHTyKh0Qo8xrOYMLRIhPh
QD4tWVGL379X/VyNorkEeqfksJFQc4sbGHN/W579u61TQ2RUyi+c/TV/oMUMOkC5
k7tXILhWoH7H6IScw1LxkqYmDu45zJYyeCPebSNiW1QxywHchlaJ0bwr7dBbnFmi
e3JVeqE8PYQZkgW/8DwIyaBx5K9LchGTcR57fLmx2/v/4VRVKBOPGA3LHz0srS+c
GJVVTS2Mf5cAYVx+YQc4yzyVz8qIMqkYDvm5x27McBMCOTtRXC8UAfvejymig9IT
QN7X5do0ANddog4pY7PknXZwysbRsMDlgbbuI0DXm0fTV99lp0YCYaWOzAMNcd8M
wkvQL44sITj4+2osLG4C9ZfnMeG6YJKuUrQ1+T05DBycyrzkDY/iZmCb837YnI0D
2mBdyYRO44NDD8ANzXzyUAGoSfdlqtMaPGhp4eoBzCu/gBtuSmgBuYdfu3J6Z4t2
H1SsBnE5sXpuJZoygashv/+o+rBI5BhVvD1DWDcCSpLwjSGhFIh1/iSOLOm18PEk
bwo6AC0q1SOhuJCmmsGTD2EZnLvRWObOTto6x5RowAyrxmUOIaguyxIwVUttn63l
jUARPCFJdK8puhWd4ZfNHF5bSwFxkKF/MCpquk+1D9aMVPq6G03yicStkzkMef1K
/fQJbyAocZE4ilgNUJmU3Q==
`pragma protect end_protected
