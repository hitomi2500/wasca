// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B1/UdwLw2eWDqYSX/wZJvXMNtNfCegGK+hF9ZNf8RY/HeBpQl1vD75eh7ZdZ6Oc5
8YyKhglZ+HACC5JYbs4FMccZjQ8doFVYx/R5TsT4F8Ud7DiDG6aHrXp3hhcQ2S15
5g1Tj2J0R29r3AmAfR+Y0QUyxOdZsNiPgf0O5E32T2w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
EUk/fEJqWVAPbBCWuI38znJ6xrdcLyWLrasVlJXjtTSFPpXS8IDxB8U8PJpXgFXH
VE7gqos8PE8ziKk78QCQYa3j/JkXLQlBYTP+2qa3WvoNgo9US+7H9LUVr2/M7XxQ
srIlYoWoPRCOciDbztfs8vPts6xktX8Iyem3cgpXhkK7mAZQs9fNHriIlF/Bhaqw
6eeUy340cnQ36ygqRO4NS6X5bfYGEypNesSZPpOEgr2iJ6at8b28agr9I2INZf2t
3h/FoA9Fy4obXuy7lhPo3LrWTkQoEy6WZr4MEjpN6yCML/YVPmJkMwEIl598EjAb
LXt8Mr7rCpfSY7CQvNe0IloAfWPMJjvS1UnL2vyF52I9mklgew22now66vvAQk7o
/cKkkPjQNOoKHDQhn2J0iPxpHBIALaOWZqhhfrmmO9dDP7bbKESauOZtOvS2Owpb
HJSa4yOh7nkvqWrupCwHiwssYMt0mkzf8lEyJHHTbm0dJhekzDLmG9AUDsBmvJZn
iwB39SVtXtcWm+WsjPqc7Xcj93qWFiAHWr0pMjW7it/at6o5+mkuoNXyj8BurPAM
MQBiQoot7FmtvXjxQ7aOLfpl6kbGREYwbmXNZ1/HxczAaIpf5QHtZG5qMT1Hz834
yU13QZXI8n+UuAiqcCAIUdrd28hoyk02b6kKeqPwZ5J85mJHDlyj9G/baANgM3gW
6WirW/rBfsQtwnc8b8PUIK/IRgHOpWzGMKmhz6HkiDQoF3Nmnqmr59GBUDr5eywf
9KMZr5N5BGADpKJjkCKzfRZoAzjL5D9T5tGQ5SWwL4PURRex4xUGf6Lnk7a6oDfF
ysdaJuueVedHLs2Eys6OSU5cI98NwneRD/83Pde6ix4mwrQomTZNZ/CKGOmz1U2F
okFB+NaXaCAnM2rpKoVongEo5+ZHXEzs85LPyw32xON0bJpfIfv3G/5SbAKEvgzj
tqQwrl/+ZfPNpa4H/ZpjRqom2cx21uZ5g5kYOB1etS7dWWuz2ShbdAqqfiCidwX5
1hufq0HSbrrGIOV9cd7jXErmLEyrkz9Pf9fCb3k7q7inu/+F9UBs3Oo7ztK0BINV
CBSRe/xIPDsh5XdDIDX6X1WroH5X60fMYOGfY7ru8cmvNo2fOhygYtzlKpOZIUST
b8MyAnUFWJXxtd5tDOEg9TowOplaHxCcYZiYgPEy19hM4rxD2foVgD0Y812reabE
OwguV4cK62Fs7ZBNeW2hBark1YKWnOSsPKsIVdtgbsJ/QIeaWNjmhy4xQpmnrcUg
JhRkONvy8/fXTuQ39TqMzOHjTgKFDEK1fUsmwLTciaATRs86vfZRfqajnMu63JOt
sMIK0zdM5LXuJqucPTy7SSIG1ZQ8H1UVzrT2U5ghzshiSWffW6SL6SpaNmzNpP3B
3m0u7mldTl7tqUJI47FMTWO0XXlhTYiPXfSFMEj8ysMxHey4oVT2auwCq3hx7IsE
We3eULJ0BzrEnTOhnGDLn1zo5wvulF7QqboCFMAizyeUIaNt3djWOKD72Q4Pt08B
okmazJH+jfq9UN0YeVvY13JJKBBOPBsifGSkqIlnpjsuOQ1kXmvEGPBpMvzCF7Vv
2XW5fryKhwVn/ttrQtnj3pZYmlQuM1RLrTJ9LEZFWBn3v+zPbPOeZh/AdBTIHDru
GXTao+ImgwvW+kAJtM0+UCaMYu5LZq34xGVGTwvdp6qm2lJ/NU6ando9ajIAkmpg
livmTtmRUwtiP4pmZgQcj3BPg5pKnjyIViTIg7004eqXuI7eWX3LzYOGY8KW9YMB
9kC6EneXTCXh0sA/5vImCXKJlvnqDcvyYvbyev47UGydoS7n985YOIpHTy85V2Ar
Y1uUAU557WsW4Ifq4axijL5mz8/vm94ITlZMQkrSxt6I9VJheAnsSQqpP2tS8/+r
cdmtFiab1lrRtuROtDIhLFBVifXY8vAEYZIXmnvccdftzdYcVJxFv+IXb7BgRmg9
eqLqnxJjKN7ordRRaPT7RFsXl6+jmbdjVkCC9ZT/vBU0xYLqPdtsTcV0RlliLh4o
1oA96nv+j+6vHvsl8+l85E2ycl2pfSXcroBAMN7WY8tDYqDEL6r0ht7lF5k2uaVz
HpaGVSeSj8cAV/a6Sc0R8nkNvNp1BeNXaYXI5bC0xS22TEZ2ZqzSWXGwi76QvDp1
tg9ZdmtxZcaPJgpsu6Q3InLhYXpiGVw1F2GvGmmMy5JGOnRM8JjzLrZaDkrARgnR
bpRhfHEl/5B+az9qgpZ6/0GUGU8thd+hLLElO7zXKtUKyN7PJMXx14nF51cg821f
Jd981ha0HuG9nvl19apCVrXSVU6oCbe+ZhSbXul61TxuxrdyO1evTx79c+cZdNff
VEk9/3r9C1V7MaTOQF+e8FpFq8n93P0hvKKsGgW5RSRlpWUJZpozVs1DFMCXHp9G
+RtlEKCuuNpC06bIuBPF4mWAbomiB6aADtz1tMuYc94vbYokQ13VdrXVhXQrsiPG
nCoHMqzYQ+DXrf1xQbecK+58EsDuGbUdFJFosf5jdKn+eLNYevlrrWvCULz6tJxm
lRdAZ+pcMw7eazKwB3gZnud2F5qYDB0dGUgFL4Jq/8py1GF3ZqeOqU/hEWD5gq8n
ia7YeznFJi3cotUB9qfcSxLoxV8eO7pa+fnSn2MM/i98MmHUxX7Xkt2n7G6YixDt
WnwVOyQWwVIeyCIJiCdfKD3574poj5Ayaysv0h2YyIgv9MD2pP+iqeU9RchhODPg
m842aYviEA0XUcJugwiKhqzlxFgriqszCzyOcu7ryH9TWyK0lC1smS9pLCc3iJ/O
0ApwA7Zy4EFp8oIzo+o+VXuIMCXBYPv3/uL/bhWdUos9RauaLmjmi92VR54p/oR7
5++SBeumHRl5BM7nuAtsWOQuWyUkcqP4XQh8N43NxqTw0sAw3OyHES0eejhrDZbY
vRasKjn46zqWMTaBuFSz97KLSE8+pRgZB2K0j5a6Da5QWu99GIUkQbxHLx/ZrWbc
Jktwu01K91EUuEcZZjwIkuloC+2HN+xdRGxh91VyGhKJa461m+yXtoxewA92/Mms
IRHcEUvoxKa9A9TqNP3iX5RT5q+AHLDC0qI+z9ryNkK3tZNxgGni10UfCC+SoFQ3
n4ahwL63quA8wf03zdltRUcXrNx2CLmS1OHynrLEaMkjGWgOl9haRP9maNaBZhDH
FXU7y/e352jn1KmELERr8ABGd2BGwM2kuALCHhNSGRQGq1VQ7xZVnyf38dTpXmGD
GVwbpJAazozGsvuN9cMJ6rjQQvfhiFllWMGyIPFekPZjc4WysTmom4B/+hSmExq+
30UVMpdywbe8Y/3X3MesHtfWt/ll5MxUi1umKBiQDiqINAMReMYc9taHx8tRZ2xR
fdeqd26WqA1WgtSOulrzZeXv8nraZGSzssVJP8BabOZe/JLQA5sy22LrkGtHRXKE
4ohol0wapg4/KXqy5I65GM8HUrEAMzrLTdhpsZZB4Y6RYHuySLzd79nLoGOLoyhj
JO16qEHDzZiPetOYtGmvAEp+nDp3DCqbCvRf54ILVctuH0DPdyjyx7Xv6Vx3spmf
GAHYbm8e6Yr1EYygS3UjmlvXvEnL0WrF6Ag+awh/Q/pL7Xj1tlpJS0l/ozm9KoZd
JTV7Efx2f9cwErvwg7VmH1PNMaksDU8Tmq7ACbMYEkehePBlihABwUZmEa9YZBjd
/CfGYAJtx5SQYnpysTn0VVl+AspjwiqKvsMSzeWwc6VspjBaBfYZ9Z/TAhvJLXOH
anWNV2SSinDOuCha8xoVIh3VEai4NXKD0a1+xrcKO3b8JHkTp7KZzBLMWDlpxjrZ
DZGC8HdHrwDeLze/P+xVgYOB+32V/HTKRiixP2/DhpgmIglJixvQj99TwrAMg7SC
eYNRGxLnjU7sEeDSs0cseHiF018sTzGAWW2SmzH3XbLBA9JqJ0RB/Mx7BgaE1zbo
3yHjxKULLQasc2LxiFHJxWHjsgtHMxbLlUdRNqZrr+t4sYJ3VzA3+VNaRPjeBfW0
VJUnHom/5T2K4huAcl7XdRqQQV+oFr9jaXIxTsiwXsuz2V0U5c1gGm4mLyszhr7P
IZmoLt3COW8DFOeO9LWLsDgkQCOu40LEYz/5Z/DGsStPen3KHcshnhxGz/ylc12U
j0WulUtwimhgvSRpc59Jedgz1uMUUrvNpnOHZapoFwAYhtnV2PJ/8e4IGZQVeVnc
cAnNW2LeR4QwcCGWStVlD+3JGSL6DaGutr81eCUq+UiNWx7Uw1+ITI6ac9g0Pqu+
H16LyvLgRvOMb3epzAogpNhq9zfVShWo/fTk+d3p0KRiZyoeYsFb9jOMVohEf3S0
Cpcxl8NRhcccjMDPYGYR4XrNeD9wnPEZDOdBWI9yXwniXJ8WvZSM8GprDeAysuqC
TD7bXyTQg0vth3cyvamToAz2ivkq4o1Sj1ipfAkYnY2Bez+7u+3FwV0XUN97Pzo2
vbEJqY0XOqRQqugvZVhZ9cS0klT6uGSEJCQS1fnY60dMsdM2z+cuzJHLbr5uOHPa
PC7QrNnUdUS5qu/8dUcINQO6z17aoMPdccYfIvZdEmAtM9AjObiUGGlPzKvnT3OZ
L+CsJIZ7H5QqPzl0NCz1Qzn+d2n9K6fqSqgebbs/PZDV5d6CsYlCdb0ZxYN7gOwC
huu9S9AJs8C6cn7lxbjq6fGkZQCqG5sU1ymLpoHiuQUOp8IpVgiCcBZQ+eLFU7Sv
+K/lH8MNZb3JDmLkUQghecIvo/1Qr56UVFMWcMYk4N8gJJkdeHAHtRObD5VhDxn4
KKy/CRaWYjV+WFUrXWg3dx/tEag9ZtIXnF9VLzo7CXRb6YXHF0TosxPVM37VnLhD
05VJvO/zylMGLPArTl6x89wByp4WcjN6hpyC7Dr/orhzwBZJyfgjhezvO/dkvbUW
T72HxqccY2RoQiJ26tCHoB1ABk9fqDK9QX86NklDyoHBO3K1lj/ay9mzsrxn/ByQ
D1nboaYc/zcbsitmEczv7ROaZoPwpvZ+Rs8gbd+Y8m6PgyJ01HatW/3ov+qXEQhC
AE+MSb2gE/ibk/AbqIshZxEvpYbXvBEVhR6Mc3kukZiysimDMDsID05CcffcIDgA
LNfBsOgR+ebbZwSOD2CpwwqMFrtfl247mfQnhijRQzDFT3FYSv/aKxyVSd4BKU+f
YXfJQO70kimu9ygwdhtg9FwSL3DhG3Rmcq9CngQvU8ngBd8yMtOtneWt1G+PaT8D
RVIL1P73dpoaVLbNsfvqCUVZxWEO45Uy3Hzrvi2df5rsIAVHHNB6uPMzEYL7ZG33
SNjw0QBgwpHYrta2Cd42vUaQG0ZDCiz/yLkPr2+7oRnZVlkoUrQDYDVGHG2VznJJ
KMpLqD8JlRWnMXjiaXupWbjQOonXz3SqFr5SJIkB6D9mjNLs8Sn4xLZmJKMCprEu
TLsrnLGVhWI1TsAWYMTsNno9UiTWcSKf8SOXCmIeOsRNilafpgJ1F4t9dnMcndnD
UAI21q5TvUiJF2BkEciiBegNrjzZVSbfgveyJE9uv0i3b9FVmOhyaEioGj4rlWn6
cXPGOpN2YdBM9YJj4FIqNGRP4TSVZ8+JN8JPD43WCKUfNDTZv8ZLJz9jT7GemW78
TxjpI7Zms4xPR4g++TxWm2PZE8mdioCXz1+CGPsgHKhiOG+FOvXfILCzXyL9dDxt
ZlsCWPQeqrgLbVN4O8mQ2HGzlfw30OjE2L8QZIP/3vKfkIhoecL2ZtnIAH5X4dDw
o2bbEEDFCE0hagfnyim7Vu5l0N+qc8gEWSgBb9eGGtyaBZvXpFXwcpXptFkzfH6V
npQ2iNgpC6zLrzN6wcT1ykhF1xieebmnBalOZPgbgw9leWSmLiwVccBuQTmHSE4+
UKE7/5nko8/xlle5v43uJHWxU/j3lvwEmoiSnfbQBK9JM80JPStrkkE0njv6GdFx
ZmWvnBZGLfok4sQpzVlAp0WGGJug86rjFGCpaYalUumMb2qHxZpIN6XEte2bvdCY
50hurJ65NGx3ue9FUZvWlsDqF18gDAbfecaw5a1o20KjUEfbrBHyEdrk5vfy8KYS
Nke95HhoU01mhvNVSZCAjLBLluHj70SnIjyaA14OHBwVuGw7ndQ9+KHhYCZlwtxk
PqO/ctaL+uComES+YqmOhZfCKhmCK9YN3d4b3QFozKMsRkB0UTTzPG7CGRy8Psez
5rcPsCHW9ret8XmHGgP8sdw3yPw/ub56xCMTwpcabPGEzqqJi19OTV62IoV6bPYz
hr25DAFq31lGirSNOKC8ScTgB0IcN08sRAoanrZaWLQOVAUHp4I5lAFAXQncs+nA
ooXPOu7N074xglxDAg3vwuABKRhQfNaNUa2P8HVQ6umIOHjZE5DhmT5gPL0zQ/sD
wYnc10YSh62qxyYVGJRZpp5EamPbbQ/Tj5zJq4A1eE20MDz3vBdQPhGuGU8rJOmq
qQWRVn9OPLPGJpWn0s1HH7+bNkIVi75VAXg0+mzGXhC7LKqhQyk4eOvg5UfEmm9W
QXvkUicuSz6W2ZBYOn3jmvBSi94YP3isMQXIVb6kixBuUR2+OWEY2U08sn5VSR5V
UhWrED6puRpAZ12aDXj8YveuF6klQ/oqHSyjBkz9o++S/0TQcAf3swzy3QbygT/q
Ni4nkWCcqoNydqIKxMpvbv3GLpN6tDB2+ckcND0+bsumgZe+pPt6UP3tYK1i22sQ
Nrr8Zb/lUJ/wZUeKv+uA3p4BJHDcueB8hiNNLh2e70vvSx6zFSs+qf98Y+LVNZze
akU05m5XgJJiYD+97U57rJmbyPqa06ifIGbb4wSnnk6wWFzxYCtbbP6+8Vu6cmq4
s6+UB+tkAc+7rhjHqGXeKL8pWI9++n9SndfPACe6kn9ByJ5uG7oxvziqu5raU7zq
y4Zqxn6PY2uwRV2wODPXwl0fsW/psRIWpqV0aCxRMznlSWGyrYbLodbm0JUEGS3h
ID2OXx1qqb5bFfTp2MAjbGlgS1FBxNZszwXJfqlW2XpsYydDud1bc/ldWTDfFl72
14leMUu/M/qmhLkWmwu8ycG1bmIm3eRLB4UmgHnMO049B47HbGvkJzdoiyiSgHoN
PMJW8yqcq/z3Gz3etkHKv4hV2HrRAJjLvjBmyty26diF98JzfQWPHWkfKk6e8y1+
41V8U5cyD9kQyvQsEBQAd58xPENzw0f8ulE7tTGWn6RXaWmkj75QSRQF2kDsNtum
blhbJojxtJAAP+It/IGmm7Jxf8V+/gyTdwhkDu5QcfQ/v0B0CeDPXuXIMRRCDjWb
6l8RQNk0z8t31CEX5eDILhXpBMDNCb8AxgR7rvVmwQc7EeB/A+5cOblnSZrJd8tx
CMBk7aHwPj5IPWUbw1CI8y3a4+gCQeqV1M52GkYai0mbhZ9r7UdQu6h88uo9uw/T
e2p6GdE+TsKv4qw9H/CbLNDqgZy3+yd0daLybUUcb0DydOSly1Zf27hGi0+a+qrc
6ytLcKhCi5Ytal7zRcRvnrWkch0n39zJdDc2GRHty3tQMB18xMCOtABQZWDFjP8a
IARK+TLD1ESKsXfJhuZhsqWM5Mz73onR2cNRmAgXxCXRRjRIXGwxd85gGkOiuiwD
jkLkTwku7Rok9cUsrxXMgzEK8nwYxgPa2DGIK8ZAjBPiqWvU3DZJeucGaX3IVLPE
KArf01X/6AgjZBl2Um4xh/m+EWZpFbJY0T+YcfJ69l8mL0Q/PDXT8hNoQzv1uurv
/RBbz0Pb+KUQk1kb5gP5CJLlN5RcwRVFKm0uyegJ7s6somN7HZeTbU7zjke/VKWT
KypgAEf5ZlMexUoLqkHOGeI4pFAxbSMXwcunux1EOyCgH6g2hweupKSpNJKyWanE
oXnTpv724WL8WVcjkxtrNKuEEsTaEvZCsofIXK2+KJ53m3fLiI3Xt5ly7841khup
JALJ3fWfOcw2u5q8kDmNJrBybCISieKKOF5OaAVWkXL2ly9oI1vprT0uG9PJ6MBC
audL11gEoXjiJSkI1b2i2F8Nj/0picCV/V1v64rJahMr1Lm3gX60nB6jQ5UOxrPF
wUMo+X75rz5/1S3t5Hjbf4V9EsWHqQlYWdujjx151oQ2PrO95cOYdeBvmEt7+WhI
4Yr9oIfsbKP/GzTGIgNz8iAk3KuBWtWgwRox20AWxwPdsElcJFeUgCJJXnhK69j1
JVtJW4tTa3U5PeXltlGN8cxBZzr3sADtV+Cob1n+Fxkohg88W2FQUHlH09OSsshN
PqydgyjSy27yYGiPvosc+rs3ZH81sQEMXb+q4zPEfhUmZ7Qli5kjo1uilBmQQlIU
Ib3gzGoSyhPjj3FPIBdccC/ADJyw5KKKnOPy6wtKdEARo16j+UcIYndTfcACveqA
JhryIsaEqvnGGcuAAuDLmVteAEI4QVlysHtg9Eh8X3X8h53RZdEq//EaEl3y9a9H
jAXx1NA+LX3ErnDfLKn5W4M36BA8cH6m3Fmsm6dUt4tl3FhSDZ3AP6TIEJbOxizE
Rom6pClSNuCXoi1YyAgL22p5mT3et1XRqAUz2Tj2Eq1v1MBQVtgQGZcGlbOj0x2c
RAYI2nAyYc+PrVaBBzPUSKyqx3vicYh5ngLr99JquKkfLb5YbAJkFXN3R911j43F
yBi0KniOJSk/YOGD3DFB3GPi/jONTQTES8f6CTWpS6G5BueW4Bz0fNklIg+pqz/B
NnEXm6FPTuBDqfopDdKfVKIHt1kQr3S19/YLaka6GXq1m6G5FQ56TYqmfN9v1BVm
aMmm4Df8XQCfDknTvW2FJvuycGvmboABhxUICXqZ2Ua4p4wRsvDacCa8l+eKJpdG
tLdQqmkBGYoF3RG901+jdom4NlQ7cGrCTINx5IPNWYxnFpSvSj/NSLMCNkoSUvPi
DVYyzg0xb6U25Rumh/6D1ykZZscUDpPhUs+/6B9cUjXXc2CvqrWX/OkQZi5rBfD2
e1ZvUB127lLQyBqT57d3XJXDDNxWY8GetfMIjEf3fQYVRx9XJXyowiC1Zj1q5SBw
CwmROuuYSXNx5jwyx6LuKnVKTa9e9kYqCJjHIewGk3SnhIAMhesoUrUKcs7W2rOk
8EYWYfvrtjh/IPX7cul96f3yLgFlzvqbKl/CPTAJpZFSJtUz+I6b/a8CmG96vxCn
oO6VUTAs1hk6G/qhw3ENCbtxG7o2M74NHDCawsqNONr0tOTZ7MZv5ucDovDo8Gn6
Q9HwA2SgcU/LBFCb0SEGBctNHhMAS4Dfyr4ch8mkL6fJ+dOPN3XguspYwKBwBR9U
BKRbj4Uv1Ica8YgOQskCoa/GrCVEI1PoNTbLKSr9fHnFGt0yeu1MnTQ1KnzhEZHI
RUVnt+T+3aCIhhg6lCw0r527hk6QKGQbim0bkxN2zNiNK4WS1Xiq4m0JQtm7fQXZ
r+n+kKhkGy7Kya3hFMV1upGtCvYBO5psTpTtlUKZzA7nxvJ5KlTrfYi/MH7FCMm5
LpStjX/GW42ZXMsOVXn42M99f7UyGSp1NC5GDpfS99uNsV7R3FxzvtO2s9pSfrYe
CTUdUgsEAloOft8uzPLZqWTuIYG7aEc7MThIkT/k6TN2Cn1nYNpdTheiIeAIDMCs
JvDo39Q5wvl1GgSRAbqzUDUe0DMACkBd2bATR2PejGsI6XTO/cNP1Ze8IhPR0rrs
HWcb/NLjeIF4brGQ598L4ILSpw5+JdmbnWKWcekIlDZN/6wmj/QIedqXMBgpbn/E
vYheQZsEn/ei4SIuhC9wOG5OslRwDa9od993IWJnKeulsVRpzcAQOJtloGW0I5Ib
ue/yP70VTGoldgRvNQ+QrZRamwuCg5KnBfqlFd7U9mcp4+Iuh53XtdX4KGMv7ShV
Y4fA41U1kzyEhPP0lgdkxmGoADIuG/hTBzLSx99jYmksUfTs61PmCmbNGjDlSods
Vkw5xy5noMdse9q5vqTK22xf/NpdU6qezdq5nuUHv9nBcTyZNaPHb8LIgw7nwNIp
OGlIIyqnV3d/v+BuzxIi9imYbzMHzNURwqZEdgHMji0lH/4+j/8YZJlBCUrKPl02
hidkUGhCwXbH6dBBztcBDuGZsEHDixHR2K9wyrWnNdRCfjmwfD1joxd6LQJfSw8G
4nC35wC4qniibNobTe7R2gUp5ZfKYw+vPEE4audDaTII2T7EPFqPOE+Q64jTiR+y
Hg2rNyWSkLoWlFr/U4FZeEoBGm3V/jYtLtU5MMP6FL9w3sLaO7n9HoJRujLAk/ZJ
9LxtdXAQKCmND2N6m+ncBZuWtUoJZWjfuGCRYrL4hX96UU4yEvBrY32pNhud/aVe
bwTShjWlisgwQctXaBCan5wdmk7E1ZQMDXffR4Hv2P6/t6YBOct3OEHWIRhdkdDw
b+4QTiwD7QP0x+fQXN/qtmW4IfEtuw/BS/2SRpaCtWP7BfpBLbrZ83Y2H/5lHC5B
NK5WffoBFsKUFFZQ5lgnL+AdqU0PyJXC48insBNB1wd5QIdgBrO9Kd9So8eMQWw4
pwva5UxBi7rbKA338kf/MkI9koYUmyLtzycmSMGDlpd9vJe6jxVmWyrIm4OHnrf8
wsXbKwrmUyBh2rTcFG9UMJLS63Q1Nhcg9uadPfDxE6ebJXgxncZzCwu9d/R1Mq6T
Iouo88iS+WJkOVwTTkCn1gRLTuCxZ4Koy8eZwM7lvldzCUq8vIkHIXLTx8bZ/YUS
uoWEnCIYo1Z92HIqNZ2mHWHAJZOtJeaD2N1WrBqzlh3yniS3e9JizGslVC57pytq
aSLjceCN95UH5GMhkElwL2r0bpW/X8SD3Cu7BDg20dxkg7RLvRxLnq6HCcFigAL6
7B1+PSpWUvOqMHcUYWx9de2IFlZBwdP8KtaIYTjjNP2slZ9Jes8x++3t2cStVdcZ
xztUHhfS3r1TXzdSf8koJR31Y4JI6JKmkOQSXb0dFFZ20UdURIVgc1JTCDZVre7U
aAeaT3/625PYSzfFOC3tJekVBjaQ3d7ygRk6EDhJ2bOs97rdq1Qh72/ydiv/pjC0
e2Pe7UujVPxs5AvdBWFA/lj2wNF859OEaMAosNurpX/jGC/qFMREomcaDZTFqed7
PlqXOszVSsr2ctdU9ZRAB2kkSO8ZwETa2oF/Bf9aog+PA1Nun1AywIPnhojqWlvl
gIls8fSMhnEKLx1ilTsFyQ+X5QrV95myA7UtVEbrxuqypuOi51K2xvUYkiOBQTio
tsvRoOXUBKptRY0PWhhxJfZAQ3OOsLgkekhhkji1bAp07KvhCHsRWkJJoQJKIJmn
Kd6n1Yd38zTH4qSu49/X58CtkTixwCvrmbE93wrpLTSvUSLLgyk00evGwXfhjN5C
rRGzZpfLe+LDNzQWxZGto4sNtByGlLvFmtjwwVo8U3ZtLil9+DHSdMyzK80JxL6d
ggs0nmGzOVXlN3hU9VZcccpf9iDSSsbKYvt4tH55/2fasFWgS4gG5HJ7e1OYzCY4
GiKuJddrc+GgonnpcCZ2bLtPnmkfpJgp+NUm0i/3Asg3iyS0sCuj7i/HXcL/HqXG
miCEdOndTgXU6ckQYcyzjfEaW4bZKJbNPALLkz0d5KjmVfeXbPCv193bYnYaXAEl
N2FkbhxlAcjYMhRowZFBGcOq/7FxH5cSmEmehNLLxgWKgG3uT2PCgwmN/qpApp5c
ttPr7FXF79SsNiEffbDutZn5ff7JXFtWQcrsgp4zf36IKGkRypIzW4UXWtZOKEqD
TUU2Kv6wEWVHmfJvlQbzdqCkulmM+mShzK8nHwBgw0v32kWkfjBD3r599ZiRmDJa
hoA6NnFecvySMWrOQGpPO02IyIPMI7QANBTlkkgkU+T86bUeR5cL2c7DMJe40RWF
9T9vO1WPsTx31E58aw8nHCzEcVb2clCuZZbudyLt1dfH8I4Xtne6YcB+Btgxqo4R
v7lU9QtyX0GIiC1Mk/4we8eGVJ3KZ7/NRyb3p2vA+MDPbZufGrlU64YaFb6XnZoN
uMeYmYaJelGQliEdxaOBWsk7Kb0hDPRDA0+iDbOUc0dRYdgI/P+Hf+r/ZSwXXCHR
8lcmztXfFfJf52l9oGHpwTi7YwlnS2sPBily8uUY97FyaN4RtX2Nwf73TDC0K5b9
OnpZIElNIAUtkPowCk67xwis1qQrIipUL7a/+Rep8OTUzjWQJ/01fTcMfHqgExjW
csbN84qvbkUTWVmpqbu94l+6Y0P+DM9jz+ULtU4Toz8YPDqEDbnhLOQ6JyoesVCv
DHlmB9npIvve+dAWY1z1gqG01yYN64L2SjXHuok/j6tSikLmBig5ldtJIhxKDae0
AUTIC060V+s+hqw0da5koOplkO1Hzovr5Ne86mxtzlPLis0Q8gjgm1DO/RXLg4to
DVJdJM0ke5LQgzV3ElCXVHAhL//l8LrQHtKIGgfIsEW9c4PnbshKMAhRdof8eQcD
1j5pcOJwZgRpRwDmWDwxhLhzdzN6CW/PljvIK4oIZV4YefjlW3B2akxPqFHChkbv
CEMA3USYra/eDbS+jlo0vutWFYuAWa+D6ocv/rPS0ln0A89kBxxBMudo2R6chBSj
3kiYytE92E/lFuKzB7QWaVvQs6bE9wiRQOxnGW1VFSsDmDWditv3bHoypMuE3n+t
HQCZLJ4NG3Iqhw9g0WyiI6ggwa90HZWDY4/42SVcdL1zCgJd93N4Xuwjz2FQcGFT
tUC7GEGptIWjKshF7zs7qzC/u8lRTXqBkeJ4B0Ir5KreZsMMrdLHQyNKCbYEN/o+
SKDlIXD9BER058uxP/qqgToNAcGPuJHQxCpAPqX1egEzZmUOiOXdFw29XglUvN19
EnwSuylxHhOyovognb2lTu0t58TDazusSCd9WnQve8jui+9cvmlO3IASiCD9whur
XeoFxolhPFgtkI5f593cP38c5OZTNPrpO2IiiFqmxwN0D4TMehuEJYu9s8IJJNTu
aRZb79EeD4HwMgsUJn2hgvazt/IVo0ba5v5VBcmCWJfFUbf2wIZV8EYw/mEODhzk
mdC3XgaLFW4VbgWUtSFjbaq8stwUzC0aCn7utqTUS5Pp7hL+ybMiX/QahvA5Ts9x
h6co0+IiH/fWbVRsVS0Lo1+zOYbJ2JEWLp5q4W/V64mLPNsQ1GRLoKpQhIA92tYT
FVsKELB3grFa7PI0E0LMQGvFJ7W3JkiS9z9+PoECNqjtvMN3z/Gbhe48FS7D5KDU
LuG5DRMrTs1Z3OUwJ7oZv/eSnnAWAqeHtrkUGy1XhBTkCZOwjiwO10g4OW6w0G/u
ZZJfqlPOTg/ks4OGlvCw4b5CvCagn3GrjOYj6SNnvduqR0MfIF1IZMLn83f9Gi9w
Ogm6DlbNdP36nu3djoIzzUh6nnhf6jHU0xVAbAhLlJgbyChoNWCOVDLz6yklSaM+
fKOdzfb7DDqgJj/RWzqvGuipzzxMLDl3mxYwSXdFj1O6d4eXfUVBWVy53LAs5gGM
ke2peBw02nVXpKfgu1BX2XiKN+DlZcUUMQhoxccajPkP+TmI6AWT0LmP5UUOi3Cr
3PyqUo933cfv0P1hWo9zp2JxAo58vq/FeJw3G8bKuWOYzlLTHnnitEj5+uBiiOmH
Ls/RjEHCfKVCUa1SQaDShzuFKTBR9m030CmXZXpCbbMY+y/SZKAkJLr5+xgmOK9Y
ff9mOu/nKb9qdjFH/qN4yL7jStrfjhwoR57GFKc8qbMgY7cqY6InhH1fXNT2meSP
RZwf8y4Lk40MT3Q5RpMdkFlVn3wmfFcfTDRJT0Jks+fzFoakgZt7DcuH8pI2L0bM
gvrcj46IuutazDcGhpzNEPb9oLRpW1oHMBG9311M7FVTKkmQDaioC7voT+pJWY0W
td9KgiiEK7bK2PU7m00ZpNt0e0CrkRemgsn+Q+u9SgiAIWwNtfBKukMyx8rvrfkB
gU0yAgquQ0jDYR2amN0JwBxnYEFi/Jl/nHTxgCD7zWt7BFd1lFm7X0dX1jacTjui
s/0KpOlHb5fLtvg8VYEg4IY4t18vbSVT64rSSXpqXb/MSEEZ5EteURZiUWxtDshr
k76H1kTrkvOt7tl1req2dfT6D3uioItoJS2XVDr7HZ4MSLbMuVY5HkUZHgnd8r6d
waiTQMyE1qy82GouEYWGKewfJ/mlmbv1V1D4cS5vcU/rCroyX7fjGQJj0azbyFPr
dVpswemWjPUtz+JNmRleyGCEviFamBzelW7syqnT1lv5WkzvniTogP3mH24uWM1K
yl/2Dx3LqIJe6ayhgyUp9YhmmnECmjmOWPpZTtpiOpjJNtkEBvebsjirxRDBHiGq
8zW5mZnI0TuZAtCplENdJLsqUtaZOX4HOLqwzqpdH8V0x5yDqouRdXw7rD2Qn4dj
wEwnWaceZDOP5HDdM8BsY/app2Kinn+sl10W9KonrMUhtcPZ2AY+v3yWWFKkmsg7
XfV5/bDeD85l85FM4xJxHGo0ud49CFx/0c8A9S1di9ilHS9rNz+msKj2sid7NhPL
ePJymctR7tNS/absDn9PaxEciVsQ8k8G6oRiHi7KNe8trMQBDNvHofN8b19gkSIS
MqunwYxZVCNy7JUZwPkNcHKUMCF1V2up8WH9ETorK9F5vKFcNU/+uMMUCTpdjGI1
4hI8mtJr8MXW3A+LZ3wg/gNCzw+73lVrJr7rrR1KIee2xaZ/cHA7BO80+7gxdoXd
h7uGP2t42AHWJ2aUhCcabh5HrTQwRr0I3nYH5cnvu0KhYp4hXmvDLigG6HJGx7CU
DCed7mHkdtmxwrjERb2w3mI+0WZFqOWyYhMWix6iaiM+jC/iu7sDmyT9fnCmxCd8
JDCssj+ggouBS3SfP+0ltCnaAz7e/0n+5Nfsb4zTlVleaePQxw3y/3CNPyuf2zNT
DHBCNT5L4zJ/KbbFLn+gKpFqVBxttIu8+6WbsC+NKDhSOrl9d5K4V4VvF8DCQSGt
hWHQSZtw7bpf5CAa8BUtMWlskeQEyVOgWDzwLeD4Gdzdb9l0HIztGAOdqeQY1yjs
6N8n+aygh7xRVT0hCDpPHR99FYBvvLPxgKLm6H+gNrcH2uunLnzdPzMSpBn2E5yK
RPrOZE8LDGjmKXb9xxggerVusa3HJi4KTn4BsrV3RBLD66VfXqJTEWYiIlQeJgqr
I1TUm+ir4+AS5EwNCkWRWoVaYulB3tUph1k/JTPtBXHKUaRG8HAqmS/8DbLcXj6o
hcHzE6NF60aQtJULmKTBo5/fk3dbcC92E1Gzx7r3rfp7vV+1uwb0j8O5VzN86E+N
sKwbTys++j8hIQavhy48iHF6QcyE3HPZkbZR3Ll2LHZED+hgWpkFGsbQ20cD6JpW
LlGc+CMNWTB952rahoyHE9O5buM97fsBmVH0QHRi4RGeCqmzixMR7GTIf2r0uVAC
UVLRE7FTguDlDW2hcoGw487EdMUiyg6J7oQnchZwYpe6JLhmpVF2i3lNezZlwO9k
2Hv0pZDIIKi0ADBjHg6j/acVJg/7ouss1zBBHeSSfhDgPBWUfbXE6atgw8wK26oT
8VZzazxs0Q5v3nlCtky4uwXkEGMwltuyaUWQz1Mv9AmpfMgmpK7fQaTTPR4+wkiL
IvNW/fHxERJAgM8aQ49eHsQc44aOCDZsBSBwxMVkUf5FUgG3S0QQOxHbVpaMLvT5
bp/YnHlp8t14fnLBsLpuwCNMtdwHwsFmmjlJR8kCSoFTPeq5v5ygbqFi2jPGK4Y+
Nx5PoXWeiMN8n47qv7DlUo2nGHKf8DZvKhHPvHWqS2z/em0bvOeeup31cdKAhG7s
GGx2FPW+iw3AunPj+HKCyqeuUA6iBMV6Fs7fCb4fie0kEYYw8IRIaXcdGBkCrOT0
EKEu16IXI5OdJutl/yU2XCSck/N6H4CT6vQELyo/bNs0g2x5vGTsJY0/QKQfY7X8
q0C8jEVndG2NNH7X5Kz2Q4Gykxinsr7RP1b2qYx43PdubOjsVzd6Bs6k0ltLB9Hm
yQlaFQvQBTsqFGz/prWqQuZEaRgBa9n4qXzf+QXQAKypJyfBfwqvg3PIeHZpFJih
HiwkamrnG0kMcrxirTLDZ4emD6NrwZKFBv3eylRki4DonaiMkDvrP0qXfery/l6j
kL9/yPlOELXt/cWU+MKAJg0v6FB6PTTIOEBYuwIB+34iiHhozD1h4BjwCV6AUIRj
U7fgP/zX6oZ56YX3EGuAHy5JSPuCT1yLP52NjE87bHpvjCu0XWQNkDSHD2fVQ3Rn
ORfYYWZAlW++ZVHEvx0DvRJlIRva47Vk7z2TW2wv75VDDG+ZRuPo47iXrsnY0rZn
1JILt4sw18k+JWW5OSlrm+j7QEtW0mSCSQFrmVMkdMtbeI/hQ5Lbc6fXOLYQv344
Ff0ThJ8v/Dj+lOLYSc3I2TOdDy0rPguFK92oXaXYqAxneGNB6OBQ0f7fR8S9tI8j
DIXwPpzw0yeJ2E5r0kPpKetPhKzg523psd/6uLFUReZEwLOTPwfDQf80Ls/rrHIL
IYx2/3di62hZx/AZGSAqWBpcLc7kRsMc6vR0Yke/vvtHr23oKZkMGan467HPLsUy
uZiwTnGV6T0DI2KNpa2lVvGGR4dTgV4fbxURi9tlpjW3/yJ6JQM3wvtOWKBTVk82
k652QuIoHALjJrtMv90EP2xbHy8w7DTdTq8zqw8HcOM5zaidUtzWUi9mKGTsrU0x
BF4zeHcU+0Y8Sf/Wx+SH66E4btK6G4+83Gz0L8vnMUHAWiwtJ014pqerZAeF1DRi
5uBFZu8HTvM4s7921Ul+9s+orb3x5abvGgVCC0Seiv5rVyxn7ubH30PeCLW/i1Qe
9c89xRUw1Hn+mwC8DOZJgzK3CkU3FLXRx334HsDlLVuqT0rKaijjxjtvjJ1XNbd3
0QySDGZvxMjLJ09FgsbuDPeK/x13T+1vUvhJe1nae/h2bDGxWApDL9bUu6f6Z8K1
4bJKtGkwIqaqdcE+36dTU80Xj5yLjiji/WxCth+qe/cstxUzJ9fab2M6IoANa1MW
XgW90NLyehLjmQM8GS4Hex4q4fhSGqEMW1AhXhDUoAcnPCzzXnpuV/ul8uLRUoRO
yewZwqiPQH1eHJLpXX/q7V+WptOepdF6mljsE3+KbyMRCvrkw/MMrxHjWSMjDYdA
wFmvCgBDIsAampClPDdgB/khAWS/HxydcEnI9HvsF2gcsu0HUbsORPEO6bb49wHU
Fa4LlQFR3MGnDcjWuBNIK4yoTSfgIkvQicfmJt76zt4obM6kisbZbd1QXD/VimMp
cVhQbhNAxqdmGiRCObzVHRNwzfXfC8oKGN3aYg7oQP/kjHI3+2IaoT9D780w5TI3
wPyQesztx6TmQm5Urg3pxX55BLHM1CreMIPD1Etq9LnINdNdeMgaOcNQ99S0lk20
05eiacDuhV+wHNt7ztZTdiaHSiLhCvjIb5M2XevIT0NR/6OeAqBvwzDMMqUOc8jl
TF2ULySHWn+P4keJi44KrIX0Xvn3rpUooQsAOM1UxGFTdO6j9hBcoqbHOQ4QZNIZ
CgPi7o9fjuCrYbEYgElmWlaGBhy2pYUp3pP/9bYWiLNid7XDuiAlgjARjakGOiWZ
fKdNX4+EM/H42hvQELTCqQqYQhawG52rRqOOpUsDwU2y4jmDvvvLHzYVUwVmXdA+
pieRbm/S2pJnLmdM378BA5sRieYcaUkx5frHhVbwsaRinSzWhB6k5Aruoxac2wlx
RGX04NlNkTAzfC0zd4/uqpgQqiQtAXUfsSSHTUjWlJPMtzxcq9bHsKRv+WcwMVQ6
Ii0u0yqCEcn0Da8ugAnNAMG1wloUqahfYrCFmkSY/WAofauhWCmMYwRBUkn4kPDT
73XHv3F+lGkvcC6n4DJtQeHkJOmC71EYBg9SKhFrQazhtNHQeg8CE6Zp3TfYYISU
78ktZHG0dwKSxFv2tkXTAyw2KbEPJJfuLnoi9jFqAq6cw/jpSveacNTp4V1sQ/bO
+zAZb4FUY8yE1SWZcQiQyqQXFLAW5zkGodlUzsK/0BCofJZWSXtjVxHtpcQlX+gp
zUTPSAv/dCYMUwf2DLMHMUJ4zMsDy1Ef0eYTY3uH2AubJfiRatgOn5UBHiaJ1bQA
OfYUdfEgTAbY1WfBd2sBMjNPxviDsvp0Mq1+n6Al2XUR2iWoVL/xOWRYSYN0Qn+t
EmBBpKomCfn/1dUeYSN+7bF4qHAe7YECgSZZP9gMYeBrGczajzHwsY7hb+YT1O9V
KA33WdpQTIKtNkq8XW/SRW54iY2mwmRbtwDkKnxHoi1zJcJcCCNuBT/ksGjTcSt+
WkoPq7ZokDjzW/eB3aHQ3gjLO3sfPjZTQXPny0tEg5ojD6p93kSXzGoaTR2yC/NO
6udlvfaXTW2UQN85YhiMbqFgpVlQqAz5aaw1cv/0+y7o3Be1YTjR5UqeE10GTt9t
lV+G5B30aaJAfu2X5z0t7PGUkjQmo39A3I1N9zK3tpcLn0GM0ureyzRg3qrshN4i
M5pryNFIGOkYIcZunIpevIbftilp9FsG9r2Jp7qqulvrjzRx5SZtqzqaTIGpE5VW
sQ9umsdOV1l3tZXSqfXI6eTx4+Cpg87q1QdWKIppzq9kOkVsxGy5tM6DLogMlT8o
1LYZpFliGJ+siPoOR/AOoRLPxIE5QHkYorIpQYpXQfe05V78Q7ZtkZOqlxYmIsAk
6rMs7bLQ9s2Q5QbTk5P76CIhlFJvOPZUJDIw2gCrbKg6eMSpGes6fjtjb2ZwxPG1
W5DSF27Lo5wKUn8wxVTURoOGAN6O1CI6MJvmM+MpGpivmHy9nxYddFTogk/v3VG2
pOfWpd9HSaRmqgoknxg5dIZ5Abyp9CPEwRwlH5tLWr/eSIuF+1yq2tlvERvFRA6p
q7u6Hd5YIZ+io95GrvcoPRGgzuYTiX087pygUCUIoyYO+RrNWnRoZhiMRb9VV+rf
D+sbKAQOZMSFvwGx5UAXd1OLgNXWnc4KC/V4q88IwPtw3g02Q4aMi6vhPPwCrqiv
kLcZowdgcKfuMflUijx0Nn9dDcHI/0H584NKVQg+5T5ATHgzIOrfNjc/kmSLmWx/
xf6POqghTNGcwxY1ujLd/unAigy3Zfpaj1ce+i9n0qfU/pG2EGumwC8+KQk0Sete
w3D8Cchivr7Vp61L1yMTQfHBgpPnq2f4RjGSfv3AmJmPoyJ5DlS0c4N+4/+N3MfR
gOVCcDqps+fxxsUe7OFxGuqzVqkXOT9LRtVScr17ABqmJvTfMYYdNMcLPDj5+w83
ROA2rY4SgZ5dppGu12c/gsbS+GeF+64LNy/s9XlG62+29GC84VZNcnIkAJxhywa2
xX+CG/Bx8lp5bkzf/GhQ0cFxvAJ/VTNghNSxVXeqmlZ/wpaAWgyqONrB5pvig0kl
BDRwQhKbuzabTBQuZsi9o2SMkgpbMExneXSj3hIU3eYRadXRG/7axnhq4ZiWTCjM
9IyLkf1FV4vveGhe/wvzvLjUdPFBvz/QTIJibvEzftqS4kvyQu6KTwG/O0MSBhWi
50zgWaQHi5ghQwtXqFIqJDTHg19rtCiMjNY9nhXJh45WLQI7zxhIayUrMCw82YLZ
DPBuIucKrutYhGhGAJ0tlar8OA3Li9rEDJ9eK66zUmV2omK6tFcu2vrVhPjQu2gZ
CZgVxPgtKm9x48T4UnFKrmuGMWXFK3jUzfv7gB+6+cJ4FtHHlDSKVXvP5BR9boCa
S/P+DksoBS4hgLGr3+XdZNCJBx0W8vpvPqPq0yO8pkyzHWXEa6eKBPNJr3u1zUdX
sUdBCVQiWa0MA52ZuoWM9So2/uSyyy3XyfQaK45l90PWmKT2/xcAZ3jiRbzVER+6
4I31+I5L7kD+cs99QCDQzh914ucDDC5hSEwc2RM0Bh5pMGG7kS44QQcv3lHgjHnG
M4JMzdlEGFDjHT4HRHHARXaZL6NDTCFvjLtRwKNoKdzVesHCJCR9tNg2kOExTP7J
5NOQWmJZMYRG3VBBZHj7eQhDzdCueI+EEN3iNSyO5El54rvA0LFLNXDRctCrIQ9f
gry3BsNRHZfTGl6WhSqRoR7iVZDHHKT3AQEDtumpYT28tWvE5R4zvgC0wviOAjYx
QAr44MDTrPil49E9i+tXz9sKUpLGVsRoUShrDPFgcSFalBUwXze5VGF2jxuZOcuB
pAwgZnB8fPnQlb+0/rwHElryQE0yx4PynqV4c0JOD8p9MRfZ/rp/e0OTWtdWSIHC
IgtREhKKmWmq6exNqQcgcScAcspXFaSMmVb74I5b5b/eMcia5Cja90DdFWNl5zss
6K1dLnlrOUQwy3xI//BFb59DJsO6SVqfRI4cqgnoyuUcYdnW8oLDD/uzlxJ7O+V7
aLkZHA/JjrwpKW5pf+LUe9FnmcCb+tkZt+Od8A79QNiChXZpnsxi6VYY2PkGwL7n
wdR/tretr0yYkc3RgkgbzSbQ+YDaXZEkQKd5P9ysRWNehaN2tNXJXrPtPMjcps8c
aiK9iu0bBYjgsY16aHh/JWNGZDLHEavj4u613moSxcOwGUJQ1bCMKhNCM4oCV+YE
vL+QY7U8JT3KAzWeMX5d+3cqSAcgnlbC5kIgctdyuwKHzdAb75VlohstARKssTTD
AvrrIsHjnpr8rfS6ReR9bjNGlfO18c06ApVbAEOXXkIhDYT0Kja561L56fGlfg8t
UMP8dEIlC/beDqQs+4kqC0ahEAQBN3FONuq4aE7cKhZpyRzAit3MlKEDuf1WBiAD
cyhFQ2TG/2Dp/pSiqRrO1R3mPGCXtwpN33/3+6ygV1NcQ8L64lwYerYT/c3A0wky
+Zj1RY6a8TZtLVxBn+SZqvzfe3MkyjBxigF1gMNEtfFdhbGF1+25sTpyKd8LNoqy
TX1Ndii76QyTI2c9b36OsHPcC9MukUgSD0vt0bbw6UnTHXx3BGmXYNFoilt0UBd9
FFgnN/06tFMInOhlQ+HV12//44BMXHdaSKK0AUENUBGP2poet9dffFA87dKHz3Vt
rtbJGwNvT5D/+Dl9rsERq6cnJJx+WvxMoG+kx5Lvbt8QV3CxDoM7ewcYX2neFkel
HZhEdpyuMJM5xrvi2ZOpkP81MSVvG+0misj5M7yUicJWubLB4SuDTHWKuoCArpTT
BVua+IIGh4E6v+k4VluaqlhYd8rw29bb4+02lvMQR68CexI7gON1nLhW6FVudzIU
FFaRv9QmL93JMiaQNiU+hT7LbSsPNDCvlMOJX54eKBYvdW+HhM1fipKoRE5kH5/s
dExTq21lGudk9PgBkH4uUle+lsu9CWbPdDxEKBDTQDE0Fp75+wJnnHVsenXfcQ1M
RMZ1+e7PD89HudBqOK/4xMGAhSkccyjCL0RMJHb1f7zE1UBA9CeSxJ+WHQSy6Ex1
qeFugJQSGxFmVJDiNmgIAfLI6g6OCiD5+FCoDLWxLU7J8VuREGGLvlzkIOvuHwDR
0+If5K2b3EAAPFaUxtzXtLOQF5wds+MLOp6Txm0UASk63g9vFP554OeaXZabwbR5
kuPIvjhtfSF3T6J/c9dsjnWuVWS9JkHOp+lz/LXPUhZmTROs4ekPYOkFjKyjP3Mz
BVHEmcl4srKje4MeQOL+9xz/K07Xm+6VhROeuHLo+VbFVdA26AhbvopnRND7O5m8
T6qNyMq9aBieYKZEPYJPvOjkOS2BjJ6rh+M8p0cN0QL0cX27eQpIPg4YiA0rybIa
tNjl9w0lqEmprCAHNSHlCbQAp7mUjSZlJ+qbVmr5p/XhcWqjOgESw7XMdlvkOllp
suqMeXTzwvUR1eCar/MSLi62WhioaQxRFuprBv+DK2lCAfqSDwIkNJmKfNuI+m0i
MMzOxvVjqaqdhuRjADjw7chhMv4ip2reBmuZWfOuOjSGHMXMjJzC30fiZy7J7ikF
dyw+NbN7Bii8YQHlkuP8HLKWfswxQv3+xHThi7YH7SZY5XGp+0ITsyeELEbkwXc7
WhPO7olqHCBNUrunwvweM79Zb6JJTJ4u/vi9a5+2iQUSarbLrOo8ZwWaFueDuS2a
n8P8YOaDuEjacSBDK8XTVG2L3Ne1Loy7AmDxWJcO1/NXMYXCTWNRdes1xuicA0Wd
xzpwSdKHThcbSL8T2AE1xU9cwdxKAxufTKy4/JrLv/XpW3RHS5waKAnL8ZWrbnVE
TPGe2CmWNCVXk60XkKAq5OmYMRa1iNzK08BJF1Z8zHggyQBiqr7wyQn7MKkQuUoB
Qe63W4/RI4gppdq+LitBr3ydcc2xODdAMizcO/Vy+ARKA8d1po1O81Hs5EKsjcFe
YjcMNK+T722Sq/RzimEdycaoqYq+BdH/DGVrf3Wl7CcKXIqEkq7rL5NTiFsb79WD
+9hATAbsAdcgFygWkWfwQVVyHYFHzO1J3UzmZUqC1W9iJv7E/XRbF7YP+RYgwRcn
dmiiqgk2q6Q9/Uhy8nlN0UZx/G+a2H3ERG9B7VYijkTVA+3GtDHrVsRJqAL9T6fK
XQN/jin2NXb6niim2cwQfHtkV/gWLWe1qb2lvwkk8hth49dFCfMb5qJWr+Bm94Y0
wHh6RDuHqnHSmLGrP6spWSxHLvnpg/mIlE8ULzkTNfiS3DMfCUH0y6qpRLk1ePAh
MA9RM5IN766GdDdxKvlizEjg/z5pmNdDZu95QS4cd3GJlcy8WqdiypH+HZgPDkCp
VrxiCLrTwzTA+DFMJLb/KXe7sJwVNPlPkFfSmdRLEJp3CdV4Hz+UanMbD33iCt9n
19YokCFpa0Oyx/9ygRegyncTl9A9GSbjGFct4ZoS9yot7VS/5JD+1rqiID+7dlZA
nL3fXh5mHpNtwRqcweLFHOhXaiFzta0jGv6OfJLdZeMNU0pwYKkqjD4QVWZCLWpw
n34Tmq67Gmi3Id7IF3ZWUvaQX32AcnQJI4nOgbeLSvTUSb5CqGMkFQrcBwskGQOX
4YQhLfgkdFCbbNEiTiaPipS/Ac+sKVA9DozaGM4K8s5GZmVZNDBXA/4myNeJfe9S
E9IANSwrp44WR2iai7l14z0ArK/zj3bCLxllhil5fCqBWoJjiHM3j6opFv+wFfUM
vU5ouCfpWthhO2hP1/+0LgoIrq6byZbwVJsRbmWvC2dYDYPzLTmrT3bykJ/zYl4u
OjyHWSgILL0SjTO/22eA1tOyUGHqMpM8fbdE0dYsAbu5GoxzWDKV7+mmbLdU3fG5
m5Sml/AbbcGc5Ziggy019R7kBjdN+RE6MAaOYigCx06wjX3RCZSn9fiq3MpkVLQp
VG3oAcC3HAI0NzrGu6sYlX7fyc66QVRKmqtw3YhvqVn0HCiE6fPa2LnbzsGK2E9H
6g0RSkVEslHhN3Q/Ckuf4UFyXE1/VF0e60hnv8KX7agqufE4XGZNhTNNC3TJ3AYh
Y3WvdqBgYb4OO48zMXdafet+S10zkQywu7eKUuvKlYJUStW3PCdaFwuVBZBBQd7B
XfvPYcw37c0rsa5tJot+Pe7Z2KOTnkIPZzJn4ZmFqOHcAK+utxo8D4yK2azTdqWV
GBVw2+vgrbUIIV1Z7L5aihe5oycJCMS/mlcvp48m7wrm5OIzopLXzQZxuI8jZQ3W
l2r0RAyi6K3pUMP677KmzicuRhPjbsbxABd/fFr1gu+ItiHfFfK4OwhKIMoEjYyN
Dp/vzXJ26bev7B2n5QVmcbwE1EXbqzsOxATELh5VN2d4MDJO7skswrqHgSTE6xnc
IUryQTgYbMrWXRYWX7+bL5lVHqoLrjU0zhUsJROWCS4Su0v/0tW2AhDorTLzt0VE
0+xs2C15vE0v4ieH+PTw6UeJpgK1SdfZqu9pG91ijgVXZh6rvBQT/S2VCDZ55atH
gSqT1waZ7UDkhLk9QtsrgKV0Hp9Lv4yuv+nqgCtYMv/L9DDDBkwwfr23ywan3HCl
PuajTB32pVaG+YOwY0qtd5wM2F2SZ1Wiwym0Aj7MCWh05vDGZCgP9pWIXzF00boI
BkIy3aKA3HN4/HpbaVkfsH5asyhCyJlok2H9q8UVix/4F/DgVG1H0OXZI06xyHcG
BCDJwh5ub89CvV3SLbkPmeUTxoco+cei8WDUm8Ghc+Cm6ovfzm/yTDauL7xHQLQ2
0YXKzXh+G8FKI/U3RQANCX5uJWoGvUy5Ne6TdlWPut6Fkj2bbwoHNzMPXSNzcQ3s
jc5arIEXryXwXBt2p8pVlttkhlIdetpp56qu2WqfpVS8JDXsJcKqe737pu7J8/XW
MnWuYevNw2z6/HdvkGxODLd8hAunymKymeP/u941BmHrupf8Qa0Y/1zQILJCw/bI
ZayjRKt/ArElddyZNINRt3U0j3Miu2yFrvSop6aFQQZnfTqRlLWTuIClHscnGsun
55/6b5UGy9DdfR9d28KFE05YCO+G9Ta5nqtpryTFatrM9ZuPVbq3L/kVAXhG/W/G
uFZZ35FEtzb9FBxPMYKgg9S4ZkY99cBvxtq/3CA7CxHogid6gPkMvG7rzy/372/A
yBWD7PW0r52C+PyNjcRr/NO1DKghzuhDu4FpVTH7D6gC4SBxZE0S/sKlSDEhQgJx
FeTX7YBT/yvhyPCDu0sNxr4MiMUJI5VMderzrOUq9LwwtugthT1JTSXA3QzHaz5i
1L4u/cU+YEw3CLZvLBpiE7eHetFYy+XLNpG/AfOSDfgWNbssNwoqbnZtuPMUvZzI
BaIWfOCaSwYLVZuUbjAc0AOQgWCTSdXlozYl0ZsbtNL8h8/n4WKYfzzsNyoR1aK7
M7h7onfUWVwNbw5kQP/MgVIKWj2iUGDzIbpTrG/Q7gdsqq1dKa5/P7u0NOaxlj0p
tv6b+gItuxcTibyWsH/HhWX/q47iXNeBDo/Melqs6t22VMq1Uju9cZz1NBojWuXD
vnnpp22vA+HOI/PnQVEPggc7ceFwkCz1MX3JT6QIXYYPeG3S/xBMTIeLT8URQvEW
cjXKNBpeZv3dPShHX+G3xHd2UmrZFPBHeSS3tb3FNUaXippY+Y+wNiDUUf7E+gy+
lBXGi9ofc2P/dE41Xhp/UH1kow+xfYDBub88vVbFhoIsZJ68Sn25/wO6SMLN6iGL
0hqW2aKwJVENbO2+SRuwbFGw3Va2mn3t2soT4BZNAz/FXvUXrh3cdNuoR81ty/ln
K8bTLeRvYSbxOezom3xk7nKZx2KWtWm7f66CUh4W+UCqWb0iB8+p5DKTiCQ3X48G
cWAhfygOuIulAsQjnNQYy/q6pmJPiMD+pZPVOtnMf+68lIxGQQHUj3Ajf9Qv6wm8
0xlmHd7GcT+yTozl+05yN1I7sJLexqq4lL9DRrO1wrRs4+v2rxrIdiOUeC4/KxFa
OF+U+uHd0pmDH9OQGyr/KmtF556XtuAlC9IAI/UdnCgU6xrbCW6Bdlm8crPRInrv
XasLTnyjXZGLP/I4d7MOCvLK6mzOxxWa6Q7zv1OcXp43oDNiG7JjixxhYlUR3zLE
IyUqb8E3QxQVo1tVW1gEKW842SAPeiL0iV08RHIbns1WY9Ew2cbr86oOh3pCSwLx
O8Pu77YVRYh3brdtmq/tRJLsJSZlGmZxacMNU95noggZkklK4H4XeVhMKAZOwprB
xJkXSQkJTUZro7/sO+ix39iFZUKG5Mye/MYoBw6+2U0UZUAqsnWHVd2AqQlmA/ep
5bST01Lnssk2A/vAjw1nX95HT8XvnWkYXsgnw0Je5e8qWDprNxH4OROQBLRa6LoG
TmF8CXffe347Ib8nN+8cZI5v2wLnPKCIuwVyjo1mN2C+WmWRmxMQjib5QijNPdoH
OQ9lWOJ3553vVwF/wV5CT0bCP9CqcZzvXQ4l3Jh7RTSIKvvzEC/Kl8O5eyGOotps
BSCkB55sgJv1F/+NL1niraVn8QBwDQSN+lwddVyvBh9BVpNHXgcUhRNWt95dIVdT
Rp7eoMpvF3rtN0XfBfuWu8s9Dx0Sestj8s0NmfHrZRn8W8+bpyHP72LNFLaU13xm
OzOQlSLSQDZzFwhK6fYpUpzGwZuJ5xp1kgScmdNe7N3M6gQ/cTfCfNx/59R1cZvO
dEcfVKhTscTH5AdY2vxZmYBfqSCIKFIDXBMhLqCb/PcOZKslVM4zdyJnvfpVJNjM
dPOmRcqx5IQS7/FWFylr86JpAUFQL99UUU/Q1DdqCKpcS1f2zjC1TZ3NEm77h+fz
XLg2e9Bm8j4wZwsDd1ogPx0MfGtjMhWa2TQEOatkApoEQUCYGYSRGyc0B+SVL/NY
Awu9lloACoc/RUjhjqSSTUYJ88Q5jCAlaJ2+Jys5dETJFRFFa+WMqVBSpECkh84D
uzcFjJwN4D7xKz+31GOKVO8cETS/yg3MUALpGoNn/qtA8bVGuW1YTlrCFlt+eANo
PIB5fDrCJSBcrw9m7eF0+cTqgxfR9iTWnygSuP2nCxP1Fz4Fx8Q6LhBkW0BsYKo6
cbhM/bC1vLEmqniQ1/2V+RLddxrE70pL658YcgIkOypz/zfeX79AtuqhWbMYBf8n
mlvn7utHgYRPA43bfsg1TOP6nlZuUfJGOrDsVNaHC63vlPmFTK6E7sWiTbSeW6Yp
Ak78paA5qv0BAkrqJN4kxrGRjMhUvRCx2+Frp/sy3KCnfAg93+ms1zkOH6GCQfmt
Ctw8TbI4iW5Zfb7SRtPlLxMZG+nBLDVPpaPxBHKb8hKWenQyiSAzqboE7YLfoFRb
/G7qAP7yC5TW3vLulj/tCNfRuThy8rkZhc0TLAbMFZ9WnjscAVOu5RMNLEZr+e2m
AOLgk9Kfq7fkOKtN2x0KVLYdaTe4kbFiqM0Prs8202S98wzHaL4LoxQEdY/ONaSq
zK9jZfXjDsP5OfsTdl9mq8AE8hIcgZFKmqrCAziMqvX3IFGSUGezgxhI0LXqK+TG
lLBxwcYQdQXEC6ZAg9gSdkbkRhK1Kbgb4uOtiumhOFO4UEi5NDKTA76Kawp9sPDl
Y0zl0xhFqJcgcq32YPFCuVb8jbt0OPXzA0TvkzkwJLw/NPionotNvkQZuvUu9/6D
YPq4n+EPXy4qMtGSawisnCqOGNeHwmsE4FIwoYgAeakFTi4e4Wh/7unU70NNktKz
4vmXmwNapq/1SPXE1Zm9b35VrpuS1EC9SNdbG4m54I5Et23mNfGNUI1P0i+fFzR1
gOWjeRz+XBd0rTZYyOca0T6lG807V9ljgYK0PvvdEoPO2d6mHttDgMEsT3lgPR93
BX7UCPPboCKts9J5rGbK3oSqO37Ls04xgRZOR8cSXrz2+3ZtHIayucVG4pWrm+aq
eQQaAGDjakNrtIf1hAqrwUgiB+StKIEja7DSTznYOLTQn/iLI+Bpt05Ze9fg2rKT
SaIVRn/hgLdBpB70QdTLG3iJIM2OokPi44VriZayBg35ovPEdsGpT3DfL+G3PJOH
lHA2IVP1fxRoUvJiODU4My81ziA8ocfLBqAVZM8AmYj++xVzaNC75UqwMPeI5cAQ
mk+bTV5Uml4yFFFyxd2wVtbkoQRktMUaWdAzR71kSmiTScnUgfK5R33jq/WbtOjD
Ar/PghDgu72c+C6QqcoiEwv5DIjS0jiP2J9SNgX4gGhddgN+/M49wiWWExOhwS4O
On5uk3w2SZICq2vU5lGpKo1FUNU+gaB60m4lXG7Dg4dMZuYcyzyYPKW6v4PVcCl0
WsSzPB3Tn2dk7iQiGa3ReaKVThFzMbMtNUp/YqMbMdO7uFQmSewhZf+ILv4slBzT
agGALS1M/LPzx0Wde6cKTg3w2XJ5n6eWoaoBQAr21qDrTE5UQZJNhefWsAcqKu7a
/I8eI5hefEkfyY9V0JBXR+5UUVdc2NTOTHVCL1hT24Z5bTRrWn8z4qIbwSr72G2J
beB+txM7fpOTWijazhqyuL7zMvYL68aksW7npFdH7Hz1GnYUYV95hHwbbsolpTnf
sK3NUiPbkL00q/HboNi6OlKVcRV2dlLhjOl52DaRikvmphs4CdNd6lt7G8XQgF8m
pozuKWdY5Jsz2fsK/rlX9naJoSaJFEVt1XnowNyBLKujjV2jK8dRr/g9rxRIzRr0
vT4Aa/ScNaA3zJXikbKt5yhc3LVGC3iY2yXcDB72ED8Qoc5IfLrBgTWx/fL4q7Cv
JXRLxjinoRCQynmSBJlunqSiXqkM0njrraWmAwVmtOLsUV8KlvZ1+b4muMoYzs3L
de2q0IWhPfz5+QTPX+9UFyAW2MB2WP/BHTTOIpBNthJ93pXzNfiodMCotGI93GWW
W3UU1oifrdg/ZzHFyFTzsNlZ4bW93f8rEFwxMpS1Bc4e0sXeYFmtI7AXe8IusH/B
rDlXOODaWQCSkln2KE32ZgzR1J5Z/84gz+pyGm5D/24Yt0LhJbCHPv+lisInMSgl
rF3MIjYFikndPY1ROud0KllGmtKVDPSZyFtspGnCtuRnelOGuinM6P8TQeI9ssI4
3pMiKZrnxnW9Kkx4OcGdXlBf7Ki87oP8XVqDrDBJDnfBWHA+N+0p+U1eWyXY+wq0
RcMxlfXgs4fC8ue8nAaCB33PBHAFADaXMjUoI4OacL1hPyNisORzQpJ6FcN8wKS4
ZCZOLUJCct1z0Gcqon7yGEQ/MJe7FdlpmBQ7PBCvepGcJb7nWL8dvf0VhEuHeahp
6ylDqn0tpXSKXPMF80qIrcaHBDTaCKtI8AvnIMxffn+zTqye4Pr3mdwfGSL8dNCO
BFVDjWDQGZrFUtfcUWgtQiSDoZjqqJPtt/Z2kmWoRzSUxbVzROiTmzPPy+8N+LEy
YFHKqUnwmyAkAAxhAzeX2Y7VXIRV8EWHBEriA585yJlnHMk7NNpmEgfYUduCMCqU
uohKt8grRhPesvsLWLD6hwHpXrzMn1N8UwT+iyjONkHIBba/KMUfkExF3mHb/hX6
mmU5xkLqLYIcrPhIH0A231d9Q9SJdL7GmTvhRbyk7Kg1WVUDUWgaIHZhx9x6wq5H
LSzOymbj6oSz4H/VJqjhUR/tvjXsN52kxkunhA563CthTipWgVga/KCdyegeKM6C
L1B9oq7PatvMOAQ5IVTRhd5u5N8FFfDR2pP4mWZOfqArbiC+eBMoeZn/fhc1wAMX
4qajJhoe5JmkeqkNRWpzP6bHg4LDK6gsrkgTJsZ9mxHoodG/47h5YWuV2LCUSQIL
XJwvNTbWFwCaEZ+o+g6q/XM/maoGBgf5jlojcwOLa6Mk42F+ljZH+LfgybWeaTxY
L/63BLsW5zifMC5ccgssKPih01dXaA4raCrQvseIeIrJKDTykbsKdjMIu5hIUIjQ
WjELULgccUIUZZq22D/fcCIbDSfXnRiEvYdqpg89T6IkF0f29ZXUg8FlLnNbMLFD
W8Y5kBxRma5GC8iH7cLN7hU8KX+D2vihm0OMFsV/iB5K54p6W42TEoYFpGZJ3Uen
HhkT6oP5BmK6dHxh7O0B0b+a54LU+03X7vYHt1ru1COWBHe4/CXRYGtGjF0SyY56
LDG3r8cHk+XIiC0VlzPGjc41hRUMI9+13nS+PuTx3sr+9vl3iHZp0VNFigfZk62F
6pEVpZNKe774whXV8I9S07CvWHvcf2damXopaLUlpj3hSu8ZrwW7UjLZ31R2C5eF
v/yAgEsdP6zGV9iwwBCgII0KDJBcs5gWktSkwz0TJx4SZGIv5GhKX4QBvRA4ytxh
U5MPjSe3MjA0dJ6JleZ46LfCGm8LHIaIDETl9yCgTsAk4VSTNE/mtdwUE0xMxOQF
GHB0WtvndNSIu/ER2UMkVdoEOS33dRN51M4PXwUKs5w58/cvTHFO5qKhXuFi3B0r
JhomYnFvij3wG14JpaR0g6o0AXFqRt2HiQ7PrqjCpuXXg8FmFowBPla4LhVjrXZN
nce9tl2onrxHzb1OAsuCEPSQ+lpcGkXgyWDQi+HKFwZTGMCSqUNkM3KDMcKLMX0a
KqEwY1zeD5NmmX/t0DjYB1Uy0Z7C02fplJeXdQ+jt3W/m0CJt7dWW1468HkQLWRw
hBsWWSY3nJHUPakH2UUPE30VPs2ftNIxJ36TXlQuRu5ibYI8RuEb0oViE/la8PvF
tagGaleI+Km6e1qkdBe7kGz1jsyC54TMaAqXdIfJSj7jL9QpWwRPFeFUdsG8Bpu+
FGzUhtzo/WFM7vo2lBOMQ6JtfQRjKxe6rKarSXVEmWFcroY1K3QpY5ch5H6Gtq15
lOOMEaaHEyswfyalPOqcjQ6dtAR2RQ2/dCcm0g8i9+koe68XaWpzcqcpxpCUszpU
UjaHXSqB3Gyu+PMM8yaCle5KUIj5o2YVI3tYet06MgLCBKEpd46ZSd70E+PNRoTn
0DsOG6RCCzBHa+0qDgvb8mEBx7WQ01B1+CWpZQuo5JydiQ7e9x4rMcdpuOGx+n29
Gucn5RkOOhYX2wJsqrWw9g//bFFGVZQ0v2msq+Cj6oizYcs7QrEIdxoX63Cy2qak
gleByZ39WjcqsnJJ+tI1ZXkkirWztjdDTy7PKIix/SOIO4yPNGRagfrRjKmbXi8I
rtCckKE2icODvQfjRV4ibqqF+S0hqBPOo6CHlBBHuf0kp9VTxjOP70qMfjaD/eyK
jgY8t/YJW01Lon0uOFgzYECKYHP0RSxFmlEE8unI9TOnHDNHWo2E8qLxrzuA5Tj+
6skXReMWxKqJKISjepDZ+1TRD7+4LFWmUYpK4MeF1144H1mWnowrajUH/8mArmQc
EsFX8/i5XSxszDTtDWRk1uQ+N5cCZ4Z2l0sVqKv2SZ0JQMS8omPFK1PuVFzoaBF3
4i6Elx0Bpwhb++/ISA1w3guOM5rbYM2rjtEMUc2IMcExJ2hqAqWNqCd77DN50EiA
8W6mL98Mv4PAaKKieL5DoKASrkEApPNWQ9Yz/k9ewlf3Sny2MpmHnkCmOvFW7ea5
qf/h7RL04+YFIyV5ZJSoj2FBjg50w1lQwUYNQXyNopp+bUJbRoOZACaDMc2JytOz
le/LPavTasKguEjy/Z+nFx322qbMi1eXFEW7ubQBG/95HKfM/cC1D+8htJY7nAYw
OtMlQAqJPhFWIr4QF1up22LrlEXM1yicEJF9yWGNibkeGbkLEwoxa7BnpnLZ7336
r58PJFdu3oEAPw5veH1+YrDv/lnEKu0YdV0AJ4X3JxydIKmo0+amF9RgV/vRghaH
+Mzb4eOLJvHMPTc5UFF4jDKa8yoNsOD5Ppzq2shytYCoOpgNgfWQfsKRlMw3OEIH
ASITHNHWJlafsZO9EW49/uLQQBIREnfW+YU0GWjo6fAa5JrNcj4z4scFKf+ozC5w
orck/RnwgIfCyhTkpuZ3Fmgl6X14bLTmLuVmnSIHIvL+nYZqKRUYrKQlSZv8tM3T
dhFaRPn6lzFhMJT1mcTcklA6IhC03OPmY83uutLHExF59J1b1/u11BjFd23aphpw
H2FlXxBBFcGnLTxlsINAScINHEpazT2yCb2OBF0UBXR2wgiv8XHA41c0iKsn0+aB
Y2t/dvXSBFMsBzhbfuntYUqtP2OK/8+j4PkQtKYFP92+932oXG6KhIng79HXz3Lb
J0ObyO6zZzcu3uvTAHviFP/pGJcnQLdlU4QcM4qtnKmemXbPxzs9Qfek6GOie4Bh
hRq9b70f5FiODEkrez8GHP4wXKQb4bBDEf9nGc+EBSQYvHhKRbTYsXlVwtWTbRto
lu9bnumTiuDmfWyNV12hNeLtWHrDN7V0ZOU4T5CIk8X5o9Eqi4F8FyAv4mWmoi+H
xn0/1CMkvPVaw3hqbs8P2wCbC/OMKIWM2W/VinZoyUflkQKVWA87xXZEx+lIf1xf
52cC2zvu99zwm7SsEJs8JCAvlzS7UNjLYZpGzKkHsv7/19p1mgdc4ovEWZLniII6
I6hQ2ahS2PVA1CrPNmCuhpzRd8NWd7gPXELLfLQ3GQ3ZYoDT2C9TMj5Q53RcxTXy
19dDoKSHtP0+HJmy0MTKEvyvSjnZpJBjnGWEQgygDogQKWwS369mDMxhoyoxHygL
zj7Nv+CYUrxD9uR9UqrS8eUOJWoD2hRxZkQc1K4bLFyte4bsFWscOmJTXSIwn3m2
yyeeEfYSukPvmzoud7bLk50lENWFLYDB3ZOIp6N0z0rI1VuNS4vsSow+0aWgNF9J
CdU3FS5ki979e85eFJkC5ZS57HhPcDagD9WqLAilWkThg6HT+JJHNK2JCzof+Ds4
6xWrkgdMSljlXr//Zi/OEQfR0RAIlo+F4mTiujq2+qj7jG53IWrowo6+QyX0R4eN
652jOQBcmYaP9FnZpRuyshq2w+Zdi15R+2vwRoXgR7vQqb46+mNysFph8BVLMHCt
G+SOw+lJAax/Z4MjYAK1tNKVVEiDkuvV5eu/SB0sG68Gj7M0KgbPZhTSWvM9yAsZ
uuxud0tvW3GAD59goCuDB00WJW+kre71seYlB0wqrsKMCeymOzEsidbsAWZ8AJ2w
ZY2WhrLzqRxNmyYhy7KsfZA+1fDwjrudPAUT8Ktztb1M2CCfrRvPAF4bPDx4q2pV
p2PKqywGVmHhDNxmBdk8rspq8Hje6BWGFEuPBxktqGttMEp6KrIzyH9i3icws5wv
yLGQl06L+bZ8e+prwtuGi0Wl1CQVDwcJzov9EY//hOy/AAWJVErjj9ooBTKW+7rT
l0915+AtRKKR7dnramLfexOqQ2c5ERTk0r2zPAAFOXrQKc6Tjh5XdDrRXufqLD/e
vhHweVO5Jm4Z+nnnNxrKl0hI441ehc02VtexVuYkPH58KOidwcWEI3UEl5jPSPVL
bHdsTtzvEuCiT+xK61HNPYwusgOw6C5ezxW68IkSAASCebvakXmiblghzaWU6HS7
maTvBTt/OP+nJgF9uUiZoSaLUdZFJSSGvazePGvgRsTVNhy/nAoPlPrJNhNaYQTx
bQeQGvIdNEj6Q3g+qQ/Q6V0b9r3933UmeA92Z0VyCXN8d+uTIyWqJsHdaO/eTvqZ
7RihKbSciQlqJGPyyySN/dE2kbiPx4sR0rvEALOSlKGYZ54mIe60LW6NjEOlQfMk
ZI5Dv9+7HCZt2pAQzHdqNY4i5G9QPINmoO9dr48isrmBhIfwSvasN93qJOUMzfKU
aJHOEeSHW6lRSYVwTiXNiijG8vjhAAtyUgQcwl8GmYXuDFG+kxv30Lc6uHkNDDnn
VyEdvUlyh5R1bm9WknwywqeTs+yW3Ag+q/KNdTt3iX2J2A226niUiKcE4fRQDMDl
6G4VvhNbqSRcYPchCh+LXgP1EVY1CJp8M5WWrpmKSUUoDVwlebITU61VlIYV/iO/
CeruyL/Y7vNU6EuOK/r0GMZo4/Dpuj4eht3sg080ZsMWq692F72PSvC4LMzLd9J4
3I1drW5G4f/17Ubf0e1LQ82Eu8/nzIyZQRTI7LHsBJagdrqtDdvEtdZU19Bb4XAy
JQeRJPXlmv8CafMF+52rlA59tN7a1mYqQ8iJ/6OyDHu2/zD7tRkoOyzsUxwgrpM+
k9llNU8ELeOo0PBpzINU6/4wwX/sMOIS5VPjsRGTxtm/1VAFSUNNxGqs2/kwPd60
/9JqHdsbKQZDlGCACg0rB7cU9dZXSn/HKSojTObree/5VanrUZtzmMGanNVfXZr7
NXpQxeFOaPM6c8l9YQ3t5kbSGeRYyA3dmifx3TF4Gp5BJaDWBYPFmi4F7yYbJXFh
B9B8Aucm/+wniQYAD9NzmdFB5m6VdgvEx4UF+1/kTlJOcbhZk+YPqKnaFJWUnuYo
OitjTzfpSqBGTh5dCZt0e/1XhpTkvufMf0jVNz9IA3drH4vx7giTBVZmix1d94eI
ArQN3nCD0EAYFI2BM/ME1J88mGXDJL8VYbU2owjG/391SYXp7oLNEHjIJaUaBqFf
dyopcv+I9FCt9q3LXCxv/0SC/9bfgxaLjHlYabtfqg5WI9xPK113KlM9tnUtxoTl
P/kEjRZirL0xoNYSmBY59jzjzx1zKDhPZtn/WFBcTFsxuy35++cD/NoAH0/FrSYU
HnzSplcVMiFLSRJJGMVbvNxzCfXDU83jQiTxs0xExiJKvcot3YTMkkTf77A024Nc
XxA0TUZs3oEr5ik3LlhnoVzkeMkmeadJ6dFpOJdArCwFZIYjbXn6CagG944WdRO3
LBiJi4R0j7xFFOTe8tRNaxXKG7FvVshEkLDjf14TEhNNueQulLEgGs+nZmhqPg56
HX3uuQt66IWgf7WJTpVXrty9aZjcy+AXDeZHXq7fqOCtwePYwL1SErLjfK5CNF2K
toZazGAkuucHh/FuRr19hjOZiICDOsRPhmU//GVIaBVQXlZv1TpFqa8bJXy0yv2h
PZ/lt7LrwC980ZGjFxG69zhm9Y7d7NJFY0kxUyJVSDeZ5lBdCDcK3Q8Au/ANzXnu
D08l19zAkwQV/zV3pa/40yqGypm3MG2xCK4mpc820J1BhzE6g32f9zI8U+5lBBA4
tOAsZYVqTkqp0edC34K5sK1WpOgmP+BO5ACsRr3r3GnihpdkpkrERQWjGD/0aLKr
jX5HqA/isiizbHV7L4u1HxLP1cOqPZr5vj8O/fImf8P3WknQwen19ZRAD4eWzA/Z
Fd0LUu1NX2RVO7ep/6M+srAwgnVVdr8NXA793Rx7ca34gcP4BjXTX7PFHiZdThGT
8fEqvv5dERE5jTPjtRooZ0Lx5Bab4a2vVRchg7nunfpD+FIjo3B4j0M59IAPwc8G
sqMnrzd+X8JaQqfG2gu6Il8HhTi4zCoyhbQKChmZYZYTD4wTvzGKRcHW0zGvOx4M
mk8BHGIkG0+0/b/hYqQFJY7Qx6MxAc+egi93pgePnAnldyX9BZ4SuaBWYXYEf3NU
VeIh4aelbmq0TK0wtF5jTQbg3/09+5rezo9TfiXzcSo63SQiNs/mDv0hsAi/nT2p
1hnfeMQSKPuVob9eT76KQ1ui+i9p8vQZ4G0Ta4oFwsWFNPMABiRCcUvXomHIpwsx
e6R7klxRB9/KYpBEYfaIlqQFH9tyuSM8+sgRnc3LzrLNnAJk1tZevwBEi9ksUYbD
Ku6Mco9+cMY5VRPvVhXOB4fqKGuYp3ySqVe7BAN7OgnlIoI7SEMlj7luWAly+6vT
hiOWOxxJ1AVBEPXjBRbPtuoJYvfYDSTNizGembEVFngA4RzZONZ5QPbXOFm1X7UU
OSW3MluGQ4gqyT8B02K9UsWTYbeoBg0s4W74eENAWdmCvDsKgsP+9mmz3Hbgo1MK
3kkuGR5+tm+5kuctM/dR0NAZ9Kw05ezieeT7LIMOJCYErt94K6+1MExVnsgiqSr/
bkd2jBkATm5Nz2GnDwvy854AliX6lt5MEI+olp59DGZikDxPFd0SHCAbfLY2WIB0
1OuQ/4CR+GXq/jztCfZdwIhzu5TCJwmYhn+kgwZuNzt30CwW8pDT8THHHygzdfjh
wHgwvTm3rhgBjxVmvWLFTQ6qljV4jO7UTq0KOuGe6Epcjip3Rxw4Otn3l03AlQ52
12+z1Td0b0a4zHzbxnFwSNYjKQNwKk32P2OtpqMIaaKSvAHD72c4j8t+7mLW4Kzq
DDRoY0Q5X/G8lKDneCARUCLthiA0tek4gMvncv4sJfqcxoTwg2HCqupS8xfLoix+
1agTpXZE00QhckdXspeI/wn26UnRv0s6u1mkxzoCLWFung9ql4GEvO1j+3//wj5D
1TJKy3M/HcvGaRhVNmrBZS1YEgIKz3M6KlmJy7Uyv6czZZmPrCxzusKwoQW+U+6O
Up4RG2/Gdwk60pCzaQPrUAhSb3p4lavN0HA7upt+CNpeNzy1ou9pI0jKw2FgaXjo
KIaKWj7P4lIbWWzLbFSC4AM84EKh78yH6/G5FHE8j4rMJwOIoUmwF2Y24dT+PjNA
8Oc+0t+TMwCqyh637AO9cxLuNqY+GNndeRIP4ozYujiUCD+CO5xb3I+BIGmr3Cfp
6Pn2iHFgSZBziLPr/0/j/gtWvtMS0Ie9bT6VcKS7m36UTUJWhVLC8PIC6gEjFdwY
Yu4h4BcIz2uac61sD3Y4tVr+1YljbDAKla+H7HtBWySL6xO4H8n66/A8Z3Z6Rwje
eZX/lsKjSLqr1jdrUJY9cv7FQgF6mzg5l93/nxyOSu/hiMk0x+FfMR0uEyTUU1/W
tpzXXsrTznn+5yMJxk2/Q0t6TiqQJtwfFwi1n6w3MwpLMmCLMLn3WsaksCLgXlJI
uX+KrV/vGpMVOvko/pEIuv2pmK5j22sspbldFaWe2Kd1pOpVi5xlG/uzGZLPDoy3
HHBH6bEl37hHL1sn7QLJhBVe8twrmUpN4ryOP9aFrG0EO0r+VcyHduPYYCoblASc
L5xp53kPvb1kpZVxGaYoSfGYz2+QVjajeYLoUDk43hiQnMsPzU2Oyz/PCHYOUohB
DatUem1gReS5p+JjjzHdVPIrr2fgBSM9S1K15UpbMaVuw9WcB29v+6UVhvhcL1GB
qDUsodobDrZW7AmB07PNrWwIhPTIDVKu2ObW3Y/lGQNLn/H2sXLxaG+907qTlZRA
YOYv1NjpeKdS+okX5TpUi2yhNenugRPhPM0gqW2N/jvRRmSuTlGebqCqI+mSFMkb
Ti9d1VI0yZi4690FVb7So3aeu3gINJ2Pk3QNew5e5xoWDxgCacPKP43CDDJIqdIY
R2xyVgAcudP/cRfZBCHEoOSv9INV54iMGDXiB3ouVqnjhjxVIO2y0vKY8RBRGh/x
IWQSwCsbQid/lNBI0WPHTNeXzUC1g4p+gRfh7F+jSwr0MQkCAMbuCVavQ1PZRG0K
03HAza5IvvBRyNQDxlfHvgVn7b9tkZ4KQsTqRll7rs47M+l3+smumx4pO8PBmDHw
vMWHI7BlIDq/4bsQamudoDOmio1fwtZPMYhZousTMM0ZaeoSLd0ztgxUpAilYB89
sGsRanbFK+po0L5m0vuDkcfG8oUWNejqBZ+8DeOOgMSyhsqf4N8yNO9urZp/9gFk
45DeP+0J2wWMxlUwdvJtNVUPUTgZUya3Jc+6+UIo50EHgIo0tOsV1ikt5g/YcBgZ
zlw0zydS4WrjOricelGwUmkx1tZgE2SVl+SexmyjJ3/tdbWQjyK8oDJ501xfFnjh
fkBZXp8SMX4dWC7sPDwDGwMl8YFkt8/e8bK4XBr7D5E19avqVLjAowAjtaS0rp4b
OE7BMxyvMq6jV7v8tqsJGhEMSjHmlOYxQq18A4/TswzJ+9R04NYIUpRyYj9XCX5b
HYsOCuxLbjTCmQ6pWWyLuUlDWUuDs97LF8bIWHLaQVHHhv+851C6Lu5SEKVQ6YTY
5gaCdKtukikRDbbvwzTrTa4iuOLVMw8k/Y6e4pCGYZqiiABo6YvVP786Pdg23Cw5
5KwFGJZ5B5TcExMNgYEYGdaqXMGM2g6sW4SIf/dkXNgoNXZK5azz9iBKKpSVJwS3
7ru3VITOwYU7gWxWinrS35oSsio/isC+oDSbcfu7cI0R0UWLtzgrxbHXV8m6sHtx
6nSFNQeeFjt5KGrB5SBSmZ5Nw4SzHA2hS1lTG31bL+Zl0Mm9qZF/poMUXsT9Up3L
noofZF9r5y1MBljnXgvB9OSpClgNKPnyVeifX2dpcEYH3IJnzyZPPOMeEfwf0/tM
DHfBkBVB9lQ0kDPHywyx9x4HURztVQHrkuPpbhfMXP4elV3wmQ5anYIeJmbK+2yA
Y1sEHIiHW9D7Di4C8zGXHr+lV3rlZyiWpDaNhP3KfKj3LcEebSUHS1o30xEjpu0J
iyNBvnuhUqR8etylzypOXjmxzh+zbuvHxzI7xeHo7lJKPdjvhdHOmNSvr9nD8bUN
zMkmeNv4840a62Mv7Zv6eS1rI0tHCTxvYEHO8oVc98nQ08YWhnnzzYpIhj4lh0+5
33wfoxeLLYD93M0rPsMENSTTpIfOnwlGTQPyO9uDk1vPAtrSswmHfQEeKB1dMYwm
w9aC+p8JCuTwlXW3d9jnXUScQRcDGSJioMQ15hL5FfJrlNtyyPY///eajfKAqbIw
NmHseUNmEVHYnguS1TBEV8BeAVMCOH4yVHrCem14NDugaj9R/lZpR21nU7YnVOv4
y9Q1N30aCHJkLjJJ3aUkOc5BNYAL9ItLUN5q0EaFyX8OSLKaxuR4VMGb0nVF5rfE
sCgZ5LvKcEv3S1nrHe9OMiz2hFHWMSP++ZR8w9wNNFgbd4xOxSD6TxKbMykKy1jO
BIXE3Bk3YBHeAHSX/CIURlpOBaVYH/iS83w36lW3R88a2SrMdwNLlPUGLSYnAEbN
6tc4wkbn1+/tC9zGOVecTRtonSnhdVE//mEd5h1PSXAa9UEWVbCMNA4r/LH5pBam
W7DX9gFhoqSR7wziXx43Ct5//X3+7wUzltwrmJ/+O33zvQqlOL6ulFfUcd0rJF9k
9YKazoMQ19tScT8tIqazWoCkj1rVWRlMNXwhczbq+sju2aciM2H3pNvX38D1/jK6
Mg1jy8M9ImNRupXW5CL0Lwe8exxUNS0iuB0SnUjfeERAQWXv9f9qI4oFmGgmOIvL
0DlI300ZjGEXc3iO1NC0AI4+MfPhiBNlJX5r0Jb9AfubPuK29l9tZGRl0HZDspy0
Go2Im2We2+CHWS7SxEBOVEw28V1Bo3ToDSjDRGX2loFLQ3c2ieR6Nx3mVa3kIJNi
fuzCo97F/YGfRTAkUlZ+DrxeNXB+fQW4D4Kzcu1l0d+/4tgfN/LMDw/qNCpbDkpu
D8u5lt8wGzaE9Hx46PCeiS7uiMRw2LCVMnFUIixOj++BYmrRb4+K2I2KwvRFIJyw
ZGtCXFsLYTEl4CS9ksuJRG+B3SM8A7OHg6r7Ocua/IVm+wv4GXorBIRpScjlw/wJ
79JIpaCZfmRMNhjY1FkZPBl82f4VCDMV+EixDN8IYEtHJCpC24DUw8q74O/PDX0Q
uvjulpiCIe/Rqz5OtCDVOUpOcnLIrx8PW/ZxJtFAVZ/w1TCcYZYglf3NbyHOFn/g
Y6Bp381mGBgOM5nngI8ZsllcW2SvzTbTaJnXz8TfW+bF6fw7noNTAQ8MP9GsQRqN
ny7JfhqC/Y+uLBJyybvDqAHxE0PSbpDrGCZ2GJVEQgZGeavZ7yRWPYTVSOYyR7H6
kJNkjB4hTOQiPVyBJbpfOhAXkPZJ7NTRLOHCv3k4w9aNoFLKH0ID71A+rLcQ2+Jb
NyVASSuOMtTpzFVYshF34hP0mIjOTX7ICDIsj7R18aKl6ZNNbhmWq1daCrnH0ppr
0Wbr76Je2p0/N8Dcsl/E5vSfkIjejbNtwOjwYUU43kqpG9lxA+5QcH9TGMsm1L37
9Tgoji99LWsy39rlp6K5GWOGd8dh21+ZX22mIbTIQINyUNrFuHQGAuIZAqvwoHJI
JKFhF7E16VjOukY8z8yRJ8o3uv3bqs9qfWVFEeIhgUJFEuYVZM0mR3WT973hY9yp
D8izySaPh/WZ/ydEc3YdI3vrQcxiQuWSJ1+/HsGxE7OeHRVCryQQ7W1Qt50j9gNc
RFg+ge2tY0YGyXVsR/I9Z7YB3W//h5gjZmKpbsaV30pximHdiO8t4HdiYmXZUKRI
XTTcCRDeaMJbdbVLD26eVvQZPTNk7eUuwBMzmjPmAJrN90JRWW3kj3BZxxNM1XDa
hg6C1D0K8t5KV1Rei0MJScRSF8qEAfGwe7pqvckXe+zsqiX2f4QAYz5Vzsete3uI
4gRHbPXR+dJccNauGiONUZfcRJZ5Emh0ugJ9lS128o0KPn23HArpg8Xt6vojbOh8
D4jl2nvbV2HtVwFnBUEdWsersA83VL8GA9DQ+R0LmaNWgBqu+1cAJlYNrkShfew/
XSCDcQCyeU7Jhg6GlHUGZk8q3iaSFpvAPBk5dSOR0+v6wCfxEwJIvKHlAaXhwmYx
TkQIM/BtRYQiPrGfugnFbmjzHK/jI0F9YNG7P4Nl/h/3J7+bGGQhpOJfiGQK42oP
IV2jnU6gGRMdDDEsgxorV4aQgmPXaNRypEPNasB4yqiolBerfSlZzhDjsfterCdV
Z+jhzp2iP+42rT7r5hNyd4kDOto8XMBBKnI6F3Cwtji1fgXaJvOvdvW7hAEjRdM6
Kb10O7MM4DFdqIoLB/iGdFjPuK8ay1P1RY3dcCs5qOYNW+yKhx0U/5REwF11N0ui
pAy1WCzrQiuDJb+BpvVLXBKjlc4ULuybFoVKaaVhquHYzQHRE8oZoLdMITwRlJVP
Zk9uarlgYoQyDFYMcrQQaurxuLJGOjK4Y9jg2pxNTIUFOXSXFBq6LqazxwPPx6Hj
gZwzWbv/YDgGcGoU5gzAoVfUQIGhxyQsnI1QfYLpXjzpzcPZdjzMR3P4Ccw9fJQV
z48s83eQ796BHy1zrDlcZNZhY7Z2FK8PWyFAT28CittlZH+3DMg8NA7IAdXL2lBO
0IVspkVZxELuHvjhoUCX4w==
`pragma protect end_protected
