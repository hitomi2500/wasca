// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
QUNkqqSXfBrlg2n4BhN0gNvFXmSr3+cldqROgvcrP/zjInNhB/F0APIHoWiWwu5Lon6c/+/XJhmX
DwhL1RFjLvnqtncQRFpdvzam8y6wQy5cezpREjDBnkf3r/BZYUEj/ExqGSslBUi+YKEuKzOxt4et
AeV/DoUNTQM0JH0kF22GFsZlH0f0WglPnyXlmEuB9NSe+hAoe76FWR5TqGo0PDJiJ09ku/PzOA+5
fbp0qRDqLVQRkxQDr/h735qmh8nXwh83CRb/WD7h/2fRJtu2yeyTHdh3JcEjxgJQxOypHGwX9w1Y
Vp5sCzmlrX4skkYH5o6XxWNi7C9+7MUJggxSfQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
D71hhwOjL5pYEIzvf/bKEJicYmKK4hzXXdIVEJDz8spQd1ogVecGTBwrWK6HePIjOF9I5+L1NxNm
y8oC7t5R/3u61ezvJUp5DUSKQvRrHx7jPazzWGRZcAIEswiINdR2EDg3l4A1cI43VyFQ8a2jlq4Z
Ku8myOhh2yRh8UonbQnsUmcD30lwtk2kx7B5Ju4X+QJCn0TvIEbKurlxSGR3gPfOMd4mzHWV82bu
JPvhv4Nz2nNUg3ZnZ/v9O1Gf04r8dLlwwiKbIi6GPfUoqNOShbZwLqvqF+k8aDX6y0mYTUqvJ/Mk
C9z9QpLOUxswNs6IKR5kT+EopU1zlSamJn47jST/VLuVsgg26RYn1ZSPLwj7hCscF4+k8dmUW2kK
+s8R8BZlDAXkS84ZO35rFZObiUG/4KCl6Sty2qLSqikhXk6yhAwhsvWgSvYnM175nvTKMTrLeviZ
NRH2IxbD6KMPf/dT7zNFksVLMaon7VwX53KjiAOliFNR21mr2GWuDvFmh1ZZJYeIVOGTNgH9C+mM
WC5SxVTornnXMG0oh1Bv0U2cG9MwC4DS7Xrv0hohYIZGwJhCT+I+jiz99kmWZEmVHPTxskYKo2+H
XdAGxPEnzAcQf+YifUYA5zZ6oRgzS4auEC8KfpDLavpI0VWF0QH8r5ZEfeICoc8ou0GZiCsemki4
sEc8kEPkHlW8Sx1jzE8jP42Yfm0kZFTpbDrOQu0XC5f1Cay+jpPYjprH2j7c0eBkXsO1j0Y9YlyH
uWWCzV9WbK/1Cy6c8PhhBpmxU8Aq45XrjReyuU+q6WKjPppSHHZ0pieFhuiFiNcBttCzuu5Jq4HV
x9qHpxQ67CJB4rXsfg7iAXmu0LJOovBQNvmWwZcHJDc5Ol4TuqQwrA+GnQ5wotRASgeS8rqxnvCZ
cSnmFNho5Yc3dfd25dDIcFiHXxHWQVJQ94qSdUPFfZ1eRvmcwUx7zQ1K50zZ2wsZvrBDXX4mr5kH
964MdvcjUTse8NQ1pvFYj4Pb9Pwd7w5dHoUkEcwqE5UjTJfKTzlKM+Kvxi9cxvDUZpKoO5g0vllt
WUMpke5OxCAR04XlkoScjcAXHI2T34BezEZd+RzgNf0pMm/Vi2Z+wGRLj7+0GQkEKj1R78IskNbn
1KrAb5qCZzFKSWpARIWEwk53+DD5K8JbAxm+XmxfHSxLaBDUwdhWvsyWn+3HY8WA0ra/GZXHv3Vs
2lb3x1WnA6kvW+9F7DrCRvLqXGGeJsUrTB2vYFsBQSTUUnyTTlVz95Z8m3/c8EVmlMgSlQDFWWR1
b2AcupDiU31bjv5XvXS5nYVT6Valtdp4UqiVUzkumKWq+eu/ry7fHQj4MsayWnSSt5jqam4ACbeH
H26D3Au2WrmctVRz7psmJRG4KaEjlAYQxp2iAT2gYPSCO4uf6flA2q9iLNYOyIuMKs+gH7IFbfTH
M6VritTU/EhFbvDuM65Te3MIXcB3Tn6TJBRYoIOHwm8keSmsx3SENw/lpOG8FQE5UqWO9KkHUIcN
K82ludU3+BsSMHfj9TXIZATKK1HBre5Ul6OUzhMimSbbVeFHrTcXIl6T7nXAKvFrZv1YZb6ChUor
1DS9WduFAxxnjquNr5+y46ZCZn3A3PjiTOEbBZfIJNHT+LxZ3DkHIU4BeFfpIfQgLLSoOSXbx360
rmCmddPdUoILt4DnYqvalRyKG+qQdBtL02Q1P7rmkt9OaYRC2Xa/EjnD/76kmDFX+rJCwU+KHaFk
Z116xfZwFgJRsjRLnE1Ce6O7Dsbus84dJJUxGrgdO4ShJpB6l7115GgrCR4x7VerEwTXYlOseGbb
YX7+74BpLJV7fmBmiQf0eLd+n0At3J/Lp5FF+Rm2sjjoFjoSCiBt+GqN5XTjiLD5FBc4DhR3EG0O
dM5aKWSklKXnZ+rMTAj9BGCfEby7uB/kRHKG1sZWuCD+GxXDPE8WWwwjDbkysDub91ci2GN8tusV
Gkcynz0FFjWZNPEmb/9b5TogaPJgKAfX4OiHnA6G4mdwz0OlEWfS7ZP2l61tlcqqDX+CKrgU81Wz
ZP3rffLarjkHGYCSASJfV5XUuNimY+W2FqQKBo4LCIhgANruE2yvOCYobx3ANLZGEekA2xVax84/
ltdRYfuyib7hUWHqfvDJx+MfFjhW8vRkBM8pyVH3NPlFnOhRq3NhrwSFc5eIJFuD2kz0hAQBKSaD
UGPXIEoEv6iA7pqVtuVynkHGqnvOYlGaWj6uKMQyCe8m41XI+w10bwQ45f9j38JPLvkj6/RFIc2O
a4JnPshZPLlGrMlqvCsQWFZUSrQIQhGkJdBvRy1bjk/VrFyw0//88t5o1cjIjpb0x7UvqhApALjX
i8MjeV/wAYHlXqWIMODqnciWg/4wg+kcT1NMckmp5cgHUl2VO5i7MUgGQOiTjeVCP9i0xVrn8MJT
4uCrBLJLOg8lBIf1pz34y5orWqqnx0i4NNMHFxSrfkLAxE9mVqrzcMd0Z5zilIoOkqSnvrvQlZe3
oF7vgfwPhk6EHjAz4+hRNeg8/EVOHEOHae+cEipF0Ku3YGeZEgpZjRjKldjJSJA34VK6V96qtHgj
6HKH6Tx3H0pw/s8LSjvHEzeU2zBzoxZC7VkPplojlPO+Z9v8nzmtqsqethpLgw9YJ4k96SwhGweR
fA9zMDORy1DBRpsYcu3vK5G7RpoyRhoN6duxT1Ad0zk5+//B8InZ+Te2MkRu8bv1oVfFG29Qzki6
eU+PHVWkZbpeA8EtUAtDgg0vSZIqrm3WsVqCjaJvICswAm+WPcR0/g+SorIbsyieA2Yzz/b50+oc
9HDnJeGPMT/YyyNx9aNnIgUPNJ1K+u/YiOdcPp98fQnE3SbB/AfZzhEic3KRkqpOz0tJLSugJGRd
pyx7zLLDZaYjxovqDP5y3POpldereJcjw03sEos18PB7WOtwhSPRJbbsn1AyUI3teiwfJzCH/5wd
LzHGAN12zqAHWs5wBGUdRKKTE3zkx00E1vI5OudrOVcszdpZzLG+n88luSzrdZQY1bdUA60lyj90
PM9vxuUYc+6EBU/1OSYS16vXINhPV6jg7GuUzFpB+Wu06t/VGiGgUfwM847OkTPFgXhouegGNskS
VCRUWcIbErzEHykQpDVTBNpn0v9aFp6/yGajFVG/zYNa3hexGTxW72SldHBnHdDCvDYOe+Re9ScR
+Bq8wT9GHV6Q/UTvH5DXpIoupXj7EcL/GJGRPt3AmBwpcwyYm9y1cfu4PJ4nzBvY2mqP2lKpLWYo
AQsZKTjGarLeR1KDe50ahmzhc/VbMMQkLy3k9FQTN8vU5qmqFFB0IzHmXLohIrtqIt0SvEtH17k7
cXbQTMtWAOUeAe56EeBgRlC4t/+tuUudWVWR0ff6YgdRa5OTPMgBAM5spAGAfvLDre9+Ary8ZYA5
XSuXUfa/iE8aUw2yyePGAKVhubfnXrgZ8M945Xo1DOe6zmqVmZvnLN+hAlKRzvKkxX7KgCsZd74Z
f0oulWiSKGO86f9XGBLsfQWhwWQthiSnwbwyMKDIet/Tbh55CwPosR9XDFBdBBc1FSlWStvdh/AQ
J0bO9bX/RBwB2BUm1YJyAAq5VgrfsjyAx+0cf4LUvq8/Wf/N+TqsxiKODDxOZyy6Z0p9rKsgzxTk
ZkOmi3dxp3bH3uUJ5H1FfP3Kyo4HhJ5BRZjcoPckmyQqTZfwaNfhVQ/mAcL3akT1AZ5NvELvbjEa
Qf1OaEtL0lHcaZ2j6ON17boSWywSfc3PqQp6kgZRM8DNIF2RA5SHjPuuf/yOcqfeTvLHtVmeH9N8
6EYiw2trG/Ct94t80/agLsRyIR2cygSz2uCcercjqcZIHAOTBSK+8oSo7FuILMgKlpv911yshovl
oQnOT6ZvRUteVzZ2b6cWxYgXohvMzRR4uZhHZ43F/IfcyQoIixWC3bS9rd3cXB+I7l9MNdBgnzHJ
SJESskjzxvg2xfitzAcpc1mi0gP9Raxh5gmX86zilK7oY74tVf6JoeGfO0eXK5l5mszVdHJdvrkG
gF9ZrjM9kNy0a7EYiCXTqDOKxj7Lt4iDpWRYJsqS6jDzaKSwlBt8z01Iboi1dR9QUGXx30mEUiuj
1OZG2ucMpemWF2mqDVSWf+diFJF4gjuu2+8VyioVhi9giIpZjE/Zlzoe+lVZoWczxwDeZukm9ibB
5Xhl6YY7Qxg39aNygMZmQ+c3nDmj5r8QDwUiLUlNeo7bV+Pd+6S828AvLJussxpoNw4rzvknjBrK
4CihGM3W/QPAWhW/85U5PhYtFPOHd1NZrgR7nxxlUpCCEUMT2yV3O/u2WXvW4B1ouz7rhbIi+Zdb
V1sv0GtSa9ALx6j9GkOnanaXueDKvNHF2MWRY+byfC5Gop7BCk2Ait2jaVmKSpNzFiLp24Tz/c/c
CAZCz8UtswgCbk8c+uXJL7Hlw1Fid7ZMdIv++FHbEZ/N4y6vvRiftWNpK/rUderreyDuaW9dLhNd
LG3zStNtWnUhswuv6LW4aTFIhtuR8kiWn68VzfGZk8Z9pdanM3X6KgJPk4vZVumt+a65aBzVE6j4
Vq5vdMcvVtJS3CfBPCM9uM0KRgGJfOKafXHRF99Gh57vGH/iCwWLJBIXkBtnOeW+2dGhaxoB4icX
IKwsomDn+yDNnvGJErYWkCOxAQL0oYroWSrWaQUcj3v/L+5I5FJDsdeol/O3q7oJ9+LLuj/VaLO5
Q5aSJPr3RcdbJWxfMSxwulwiicYCbQLriSeorAbV1GtEh1meestpuLUVhC3t09j8FOjfN8auZbLV
HG2YIIlD4TGEWDGqMRusigZ/Y5bXbjpl85D/fcKlTJv3lo3l+4wpQdWqvj7xmNkufiy8TCukdoin
gXHSDITxhFRHiQvQG0mL4JEki+Ltmg22E/y7YdbVZgUBDuUk1uevJnk9Voye8hHQoKM0KS/Gwt92
IfCitvfF0kbj47rguvVZXHI5la9lpykKWxgypD94XFZMva6M8owXwzqLY+xsb6Sa+775jsWcQU65
FMacGkdyor6LnaycW7uxoAQAPeaMjJmeLowpGMof8Me/LaL8VTMg1xt4ijDhmCS8nCHO9p231+XE
tiX9UXLvm+FaoTmjZwYyeYFIkL9Dt6F6tlG7tgTkDDRzjC6J0tTyJTpLIxNfhrm3P3qIaJEXsa/4
kC+Q0YRrphsJ9axUTgK/Ql465ZvRFy9zLCrJES5OxgNTDR8aEFzUjE0EE+EyYLWShBzNTtUgGnxy
nmzQZtmVA7+eazi73Rbh2O5WkGAnciItgXnK0DnToULJUE1aTBTShCgpsrI6o71Hyf7rc1X2pCCM
6jOqs8ecR/ZutNDFs8ZYQF0lYdEHAsCkwlrPc3UMSPKis+KEPNwxpDtFkRWSeWFCMuZcJz2uH5pT
MtayMFSRP6INcpWR9aZPUfhCd6h9Cxz7aD7xQoe5r9nb3lWBteVEB4vzLUUpNycEzDOPiV13XAcK
jCPVtY52TX9HlaeSpDtrCJh+2JJnRdiqlAPrUsNxDHLVBJQjSpn5ZQboX6En9fmEqyssaTpEnrw9
56wvByvUW4gui7tr9e8XhlD9Nyt0Hnlm4H/A+12sI40ksnA1AAQ6ANOwXlZDCxsQ4TstGypxt0zg
gwL6LnWSMeh2PKJJWHt3K84g+IF+cMrBvHtFh1TWeTbk7HyOPCIAD+BqGQ66G5tpFMW5D0zkTY8s
k+ihUDu+DZ3YU5m7CVUuitGTac1Cyt8PebVx1hfpviGdcxFawC0XBdRIclEIXqGt8XJlPL0iKr1B
DbYBK64kbS0kR3yWh0k4N3LRe0vREB7NFXnBM2sFIdKSD1EVl6plbGQzW5CU7PzPzSrvVYlHiBU5
F/5C33Wq4q1Xrv/kfydq+kVLVzXsRWX1XzXjAuzrgpC8AGDw6ZbWwgK4Z4xxpIiJ3mNURT4G0fo6
4s/NgGnu1o6LyMdWePh/okCsjgHgyCov8izJ6mZPQy4sWwVy/NSXqmmEzsMGmZ9T+OtnTZnQFp7R
Q50pGO4YeUfk2EmXXWgKcuXviV7MdZAPle/J6TiTk3eHf2XMgkOJPJOTa4J9bRnZgfJX6ZyRFMRe
OfbloUJXNe/7WdI7XOhmU5zeHbuzAoxdLg7pR74o6Lvt2ETRXTB1wIPP5VDgn8zSLHcDAh/V7RWO
PdIBYltBZVakVBB9MJfTyV8benSyrciLmKlEAW9zkLSpTqdUJDUs8CFfs57+dbPj467L7IjFDyol
akIkcDVYFJfj0T3OUXQqPT5AnoLn5/MSvfBDIU6vRJATZcGUWbP2chQ+5Hfdu9aNHMyRhk4BB5g5
TYQTqcTX7UUWW2Nu7dxU50mdyIGpHplFz9cw9Wr0TZiHL1UcURr0ziZWHEcRalu+k0jWxBexxo97
N6IluZKzw8Q1hcXx3emm12SG88vOnYvTrh85zsn6v7e0VfRUQLnvooPAOBH5spaXjB6JrFd9hIvC
Yp+H4bmhB/Zwys1EmDdmDTBwiJPtfTKXIWo7azSNzSOj8r6xhNihbB1iP268YWExbvRuo3/x1Hxk
fh8gK42iTDLB6oxuUDQqTktcM8sXZM+SzBmanjCxmR0NRCEMMcifWm/w82fQyA5o7QDnagxtxsxj
8wCSdsbHYdqEjnESVxNHwJsOGCAFyMLw+1bCKXhlIpTjxISdCW5P/05cAIb+boVqfwVlSEPfV8yo
nBmDxmYDYG2kilZFIY7wd4NnJRwu0w7UlSUaAgQiQrdknnY1xuHnGcWcwNtjMoQFDbPyMo8nwp7C
ntopXqc05TvbH0Ukrogeo4kwywgK4lK9xuLSZBYcbW9mT6s3WgKyVtaFKspd6SFBfeBwr8qPf7NW
7KaKknFCAJakeI2Q3AAu4nRPt846zQQXj7t6ZZ9geXJf6mtpCqtzIguPImUDuZbn9f3/bBhr8M1K
v5w4EDETwR8nIshlAdC02snaVOH2KiqAoItDX8LCZOoy+zLpunX9rvK0AbxUyPSF7Tr4lGMeQG3W
PP8cRqanqCxF14m61e/2mhxPjIp0nged4d/ja1C2an4FOyvOLoGz5oUcSMu8iekLZCkNKZJeh/DD
hoSytAqNr/EiRzFbCDtvAKDwvRrujWGzR0FtcwITxgsyJGmy1QzvhqXA+noWSR//8XEI+4ax/O2V
B2qITVTPTBGmaUFjrAJtWkcJuvsNof+UzJpeC7wwMp7XWfmK/3YQ+IPJcEEa98aa1uxbNM1FLt2K
4Z2gvm7Hwd3QlsUG12+lBE3XFRkUc81r3O3KOs6AVgOjJFZqi9QLvNbIJjUN4e220fKfX1q2hCTF
tYBweDNjF+NcFmSoqzOcTzwYAniaLauA5Tt/6B3N5BkSSKHsbR/mImBgfpbsxmxKHs0rDFQZY0Kf
EZkilKlr6yp5HpZ0eqCCMEyouHsVQex9TLoSK/ktWuGzfqiyUcufvtdn7GVLjRLBXK6+kwsCrY1C
K5OB2KDjBcla+u2CRJy9hI0mnD2TsXrpB7BoIpTGxZbuHROcYwIw3Oe6kARxRxq0a+LuCjecep7G
JyhFyEFVoIEui6bzl5X2PboUbdv7tb8ZlPSYUty9PJbbG08Tob7tcJNNeQEBhOoxuUWU5M78wmW8
OqAD0Yd+8h4j/amzs73qbf3IoowxByGNL3zfEZqWAmG368QrGpwh/ZpJiMaA3BSMYGf3MyShNnl/
ABs0ZrPU4Oybf74ZpRFqzurWMDU6Hx5UEW2e9kLbjYakl7snPLq2y2QG3/Jj+6pBN42oXVLTJdvM
BmYj5t98nvhydsfVT4dXamzg+qSPN3wIiHdRf1uO1bg9uGZlftzyH3uvEGdGzQyMPLlWDcti/EZf
eJYb1engdl11VaGaew/CfF871f1tck7CfWCO0Q29sYB+yQ0r3JA+7MNGhdUnpXVbd6Qr2yoUDfB9
J/03200m7/Y3btm5JnaM87EjWAArvVVKWyY5A2Kj384V592367pzw5HE6IAqI+/i/cmWEcmSIN8d
MREzvTHexTp6NiZUL3GN6Pzfe/Alf+pmqiJCTJgQyFD9NTxT40iFq6+yQC6EBbxHOajvvZ8hkihV
JLjbu443H99cwTWTiS21HhIndcc66fFgQTraxznns/PHmtxLkFCjPMZimQkXqY/sRrw+l7E2/O1e
c6v4bNy8XVV8Q4np1DVOyENvm62nhoFmT/Q8lFiT/GrdsP6x3oQTOm3ZQbA9UycNWzZiqYRgatCx
wol62hDZheK4aKXXruGra+jgkEuw89gA4iodGXGFsdNGP1CYRHWGJDzaE8XgSKVwee3+XNGm7DOB
4cm/mrCSbO25qbG97L19Hji0brX3iIFbXyJyNVUp9d1Z8CRX5elHtoN5fZTwCf6z49Z8Z1wyQm7M
WrgEtYcDbu/kRGCZ3sJ9QQA5kE9g+oFvuvI7fVUAXioX4Qjo5yejrLlHFI3WW7zR1dk12xzZTNxK
30bTGq1Pxj9MsbIVva6XfYGU17Mj52aF+neODE2vNFg8CkCtM9KJHC67udz1l7PAGAgEwUsc3jNw
lcle/UORYoU2WcLGBjpwnV9g5wnjgY8M0ceW7iBjLxfnfvywxv/K2rztp5Cq0hymQLIulN0mWsp+
PQ1DEqw02aT9KI8VuVWIO2ZiWCXEdlVqoTTZXUn2yABt2yD81LBDegmj4xmhoR2corRcqiMG0J/U
XZi3oyEkzcqFurwe9ya/88gm+55a1qcd5Scu24vM1zhOADYJjKRZZreoEYMywqpHrKCIM0z6isvZ
EENPbEFZLgdb4297LRobxJjKTw8Pw3Nh/q9xJSLjpORMLAwNwubH1I/mwbCf1JY3vETgtRPLb4AW
3XCY97asVhpSywKs3sSYq0ALIeqD7Da3t78fJOGo9RG8nUd67ngRu6Nu2g+R4VZ840rYLMJ3oCdv
6/rmAUs4a1qxciZx0HnKjEVgU0yjpeyFjWl/wUlKuyODvNlic7wsKisnIZ20+QWIQvtuyRHTkP2Y
u0g4fR1MGIyu9gQy100q6G33ulIDfgbdMOrG6EwJttvmTzvg3MuvZNOkrCpucxLwBn8lKaTDn3RU
xACe5HS3JduKKYlkMkIQhKijpeUuXWPo+VvV2UNvglWLgGzPnqxQmeS7sKI7LIlxWZcXH3KrNqa2
adrZLx4ySgoDFwalGJ2Qq8JaJaJFkTlomMnJjPupKrZe3g2ofEEUwPXJqdsggUdRoEEG8g5Xu3Gl
HGtlpqJuNPVGCuaHwAzKYDOoXS3N/l1kkp1pKPjnIIGCLnmNPyGAO5+LJOeTjN08GBaUFZC6T6Qe
nL/ovo8vsf3D4Q5q8pbKeg9EIumIUO4OZJCtc5GVl5ETxPnUUvOwixvJeFjmX30ug7I7KJ5SwNpQ
hNcR61stSZ/Vn2aWWiFtn72AmLI6BBjBenQb8Cgl82Ap+KTcHObulHHTDOM7lBVGP4sCIvUjCGkx
yfnHXmv2W7DJ+38kuwmyf3M0FVWL1NfFPTq7cZAJqLRz09iROAPZ5wNvDXwjBJn26905bpXzvH0F
DqUysb+B+RwLpQglgcygOztkcGE7ggObM92LWTOJBiQO9PyM34Xn1ZI+nTnxsac6+tc5+deftATN
+/allEg46J0NAWjlPmhlPFp0VVTdZe5TrNtmKRuB2PM92u71LcIO65VTZ/nPfYdgKviWY4bDzKoG
c90FkfbBuDMzDBZ2XjQfZFRamuIveU+eiImGaBlknu/G+OgVu8nNUhfJGXz23UM9Io6arOld3cBz
3+9axQjJOtAHGitfKvwnZw1oGJa3QJzyla4xMnkk+JYJMiBSl/m1qphZd37LS86K65r5GnYCwNPI
AaYS4THFOf5CRpUZC+NvRkdWqwFGIj+i3ojy8mn/vHf7tstm61rRJSwVygCJBMCVkTuzUkSm2+5w
C9wtJY8GRM3LPLLxl8q6j/YkY88vLKhZNG0oUKUNRD7QfKW+tfEVTEfY6Pz1vLPU5kAuEdD+AX52
ok/rWA6D3i35TMn/XiFMdXqbJy6KUdyGZKTXRtMn/zWDwkQcCYX5e0qx3WWs0T5XffRrZAHg4NZ9
EgyeH7zvfWOeY9CHFqH0RmIFKBbL4lgHxiR6ShLdEeAwZ75G3OagOTmaAGRAnB+NOF6/gQqh1kWz
fvRJa2UWvW9NV0SSSmgXcdyIFzv377ZDpsTQ3xya/1wqxZS3A9SbeUwetJn1A9QZGYYujZ/5ksC8
7nlpgMvwa+OC22STuXfLGzjaLz9mykzhCrU4rdtzNT23zmDdZXfpIBk4jYhEmS4BjHpd144IV0Bk
CaOt1WZVx+No4Ztloj8pfbz/BqF4CqN1Xsh+DLa+k6jNp8PVZc637f7JZahT3vL4rs2ux/R7RVTj
Q0Zfd1EfDLn0YlL3mqj3jjLmE/LqoDCBEIP7xg1o/GRqihrl0okrE0iznh5l/K605cQyoNvT89Bw
R8Tc3RjDFBKRF99sMo7XOXlxbBwULBK3HR3SW0yVGeTpJjCzFPJ0HsbXDKgdMo2EVnsCTKZvGEBi
mj5cbBIeReJg/KQ0Y64pNL8qATWz4P8AlEhJFAYu0MWsxtxXYcPmlRkdUhCvhgqL2FhChIxgQNot
JZ7zKIMIDH0xRBfQ1PoaixVQCmoa2gLwVNxqqNEfL3BNb1od105FdEga+BqYIcco7uXdzxUehbfo
RkLD0nNPRtbUHhhUWiZLhehyXYRQkRJIsVwWntkzDEfmPPIwqvZ3zzM0yvCa2MVLmOkxq/GBP3UT
YKFuO/pUj0OIUD5xBPREVEimU1D4FXz/NhA2mUgi8iu3/UqlqxJ0j0QgzIiCqW6xkGeJvXvOfJuf
svXi0sCGcrSjZTnF/uWk1Zq3Zda3GKujJM6nHzqOaXTTIGmHtuSeeHuHweFupOj5AqJb+8Vkebs7
M3rAsoIIpFhFFlnb+2aqSc74RhzciPd4irS1nBQyfwQFH+sOfn7xTDN/RmOHfC7uhF44og1o76i3
InhHUVcNJm1M8ObfRtTA7K6qNHD0pVXHjqVNmOlGzo667adVbuhgrb5c01Cg7gXuC78qP38iWVqM
SynNbyeMgQpVbQm4yujRD/T24slO9jrkNFeCha4EomkVpYA928EpEhZoOAVjrksiXb0AM0LKAeku
9NR7KZCtz4fvCQ7sS5/NPOGw0aPQdSApgiNilJ5vnyu/4lAhn6A8l9bdHxc4ptbSO0fFJlGmueit
eAObXnS1MpFcPdHbM+pgo2hJr1vmuXhfORBUsnTVAw+FJhQHVNwSXEK3bXRsgwCkl+RSC8P0jT4g
eEUegzgjHnhnyg8BwRdkF30pCrksXg1KW+PDw3tnYFdia5/xco2UvFYt5nyGYLK+QJrsqnXaViiY
j/DRB7iVg+OVo8FqBAKMQcLcJzxs3zKFdxgGa/iwlbdYGKTScqsFHeiHJhHxgCppJsbNVQCKfOCs
/uts32DSX1BrfbjKLyrK1KYDOOSnhBpz9T0s1r8ZAp1AD3W0h6EgxrJdP/onNiJ1h5SzxJtyRtLN
FGFMd2vkiBPs5eC4C7dqpm18WLsRex2BDkMSm4EAjHhBSEsuNXhcHLYU7rdTbWup0h4M3QJqmptj
7CMuY47fweKzJD3y7mdzrKUqJ0oyrLRBpps2mQN3C2UPoEVPP4Uv+eqcTjuGhQ4dE/UnxG98aA6H
GzhdY11ny+lgeRsbUssexWOOUzlyIMnIaF+rCizlTVvg1sp+kj6cJ0LnaJJgJIQZrdP8EDjU9eWm
Dnj4HuBUDDI9Bi2mNilDMZTwLOpnGP2Z3f2beTs3XSCYvw6Nao/0MAZY6tW9v6ZUwdVWVzdTt6BC
EpogABrDSKdqC8mJnaVUTmBnLgAOpDmQ1K9FA8HJMzhJZ2gbtkD6F19uquqWfJ1YAvjDJ9tgTXWZ
aWkqaXHl26V8+G+6N94VS6BAi77hdoCcziyd7qHa0ekymqH5gKH15EHxDFhvEZhfbOm8F8yY1WS7
jIHreXIwPlWt68OD1B+rnqUwyzPUjZ9fMTECHWIenkw9zLohgCdB/9dkmH0p0tyJm+DUw8xYIFea
Raa79v6rT4vEEDEFCW6jMqYmGhxRmMnPjoStw06LR+i934JfIrnXcctFRCXDTvVmT5NUh56AH0tr
QsX7q5eLxMEgnfocoW5rkUnAyJWED0f9DYUm/ZqUO3i0Vmqk11hvaV87ry25mlZGRidKx1/IcLCb
aBKJvuJCHCEii20l0s/pojeyzm/z818VyoSE13B/LHLEcRt5MlsFeG0vvaR6WqE5QFeyDuf+29nZ
7UL6QkzFu6US/of13J/plICXuGqj/d2dtYrHeaky9uucSJlrzUjJACC2pBBHIB6qiQbiWxlTlTwJ
ViY2UiJFZScejo/DLwR9fNfUdCTsvKAEcxdBxGGhwtFhEN+pwp1+Hx3da29ODA8PxDXxRtOizlcJ
+9N6nQ+uzX1ITnwI8poZR8/t8oedc/xBB2kvHL/gDcML9gs5Zk2xbqGbl4Zgx4hir+rDzJDKVtXI
wiimWx1ElQakaI+3pK2+wtNVmtnxMmBvj9sLSMzHLhwmV+48HvM2c7l5cadMJt8wM6cSFjgDWuo7
1pMhuAqlz+JH3Ly9rTOUyHfLh1hIkQ41bxnj5xE2U8dcF7KHca073jFOog0J8fRlVEDGLS1maVox
RdYUtJ7396G3NIbfBBn8JOqG4JCebdXvS/31E1ObVvV6tOddrMaJR31Wa14y9BmOpg+EFYQqX4nf
1P8IIP4joCDXMWj6T76qAOeRt4YTQsh4dV5Uw97GUmzgKvyFWvLa2N3xPVTwr9nBhUrjT6H3zzYk
e/x0z0fNulOT/TR7j7zLuzTNe75N82GoFV52BiL559c2MvzNJR4f8ZgFJM3ibrsD1ck3wognqu28
ld02kbPSzmc4BKurFtTVYpIjSPgQ0741N53h6oRx2S5cJkc2Z3WSzBI9Nrq5GtYlrnonjmawWQSj
aU2xPwMmwF8UgyEFyikBP6O9vGIGsAKretM8etPWORx66N/7EBHq1CNLr7PYLwpSWIxuEJBO0bq2
7fiKf1N1jXjK+nUh5XpBlqDMlzCPUSPk4YZ62siVDpZ8tyRMO3nNolHEuQPVd83YpRM+EwwnT+O6
GfXx0e9FmO14B8Bpq43r8XtPVeT9yQ31GiBkWjL/BPRJDih9QCJpFbWAnZwgB7Y+EiQBk9vQUql4
Sni6Us3RXhMT6YXbzZ+t/kQxLGnd7ktLXUvwa6wPtWDMdI4banGMDpvelSklO77Ai5BRkjIFjHnC
EE6zGh1rZrtSkyvu57IYl+7KY+82o2ny3CwvSxgO1GEbK88bzeAhKT22tp9ypIogso5ABfc1ApDk
5JGiJgPTFKTj64gOTdKEikIMMAYUV7sVptDYz9+mP42WmDA380XXkZaxUyfroSDseL5RqBwZD9t2
aqC2EUaQBpqmJgTKr+rrLPnKmK2+vTslSMnslmbCAu8JlnTyOUsrfQm6gMirvOtegPD9fiUDBuYe
1yZMk02RoYBOkCb5mYYe+iCZL+ZpXHoj2mGRNK6iiKPTDzUbqfT74nQ2pJTNiFX81Xmj5ZgPauZ0
Ra7rQbRtdZwcfiPuQ8aIfe7oPMuYX/zdDzVfmyF/1PCATF5FTjuPRxVClz+BZjBE80H0yHbFsb7F
VwNm+CIeFfFhElGySP4505qWGuZElHQNouLMIs9oOFDK5uEYhC4G5sU+CcaJ1ImvpQkXWrWST/my
VuP99Cx+UgJkx3TmTReIceFDACUr8Iy+MeER+11aNVKD67a2uoUksFZapgXzyyDNXT1V65iswssx
S/J+QZDTzHbOr6YJC8RNsyTxrebLLS3VUaY4n0lXK6yKBh/CMAmWvBb/dLzB5JGa9AV4ubz7CCG1
XVXfhGJmHY3lXhZ+aZkvvNRltpL33bmjDbUOas+0Zz309i6NZLkDWcCRXURuTaEKJYt01JFLbnc6
rhQxhBrnS1EZoMbhIYRy7Y51lG17yOWG4/77+ePMIhvyyRxg6nNpbYbwFpKQQbsp4pxem2dJZSW2
PXJFxI+PcCJX/UJ3JQhWe2yvc9tocqf9rQEyEOhu1F2DsTuiS76sfe1AQz3zcAwNemwuZmIGzC0z
thTUsKN7Y/LMiuHh29hvFVSyQxKMCPawr+3qvgfmmJoG6nJv/QPBCcJDziW3TT6LaQ3IZV6zLtPd
l0VMz9RrN8GC42VABdFrriHSBFk94Hg3kSA8bltaumRTb9DqIJfSItv2aXyEm0qfd7VSi2Ks3yFo
zVR1xq1KfG6tlF1H6JSoKQeheaRa/YczERulh9LQaPkPrZJ4SHXnElqOqZe8rZB02Iafhp6djvuf
hEGOHERPQ+z0QL6nCn++O4tVnj8NRMOkJ/7mXQrZVxuhjUIIXru3eISnz17ZeKlFRJO4NJwrUVO3
OH4purcRQVfTUMFsQ5xjfxcEAw+MjlPKHdX7FAWKWeabaxiaA/iP3vy6ctpMBTf4paz1mhRxhmIS
fPjVK3FbMSwQVgAwVX54dwd431nNj/4wJrKLKEUyvrJoLLADUERzPugPCKlY/OgrMXer9FinEXRU
NfIkOR194NxXEwcYv+KTUNHhoACmIKJsf01vq65dmy4tkfhL4lGEy54Us7KTZ7pZWLpeKPtzUk9d
wupE/w3Ly0S4I0ytUsVTK4lk32/3Tx06cmjiOSttx1xpPfHyoTAZjBa0DsssSBgKK+e+eHqGQIF8
+VFCvuYA/yFRJ+HoJVeJxJmmbFl4y76LNcfJMoCFdcG+1FHVljUQRGWc122kN2BnBnKwUtVx4JUU
rc2iakXONf+mzS4cbETxtSQv2/TnEzz5RA6SD2MsQVEQxRPIptrHE9vPixZAyYCvjOzOP9PzM5av
4lgE1YcEnEBJbTVRjDdqHMqUGeirvWwF9I312lebmzQCR7c25LvenJgWRbtHja2ofNJW1VuRNgGK
FP8AYeU2IwsXPtw/TX+jZVJmFdJhwbJgTbnbP1a7idgQKS88E5ZxHj9nSgqOlD5ONUwjZ/1LkYqc
I7mFZLoiBO3KMlCeTdgUy04BY3F8El9Fc3Zup+wga09A5Gy4au1RVN0xYGdqm7055G59NC2/BEa4
3IY8CMHDqVqk4lSvBb6Qzx0txHmIpI+k++Uxj9UlrJ6B9r/fqp67Y/jU+PjdoG7Xv3aM0CGLfWt/
IuYMtHRuVut+l8agXBY2gtCuq96TEG9y5XRd68sb6l765PCn6Tcwb5Bp+g6uZhQmRBccYhq+BOVx
NKuSPZDKE0jZf/WtwRbHpCnQTZsQ86vMucRbLhDOUS9dwcnQCKmPOCx3EJLxRUCDL9WoQ0ALC4if
C6O6PPNo1csrZY4AWa9fdPqpgVLtq+1S0Dv6a4JCBpzN7tJ0MA8Q6PDpkDx/fzGRf9Uqnw9+j7Zu
DKkYF0wApJ+dM3+eiEY+nd2O0KYfXFW3alI4/Zv+dfX9X4xrgAV7kxJfbLOoL+KkDe0/LQqDU3xO
qWCgxsj840F9m1qXXtqu3/iQud/B5+4TrnQYNtzn3whcaO5jFUQ6eg7zHDEuKCQnl8ZztfHtREBY
T/sVtDrnV3zTp9CdPiH6uF2yb6roCRCGRGYXpP5sNnUl/uVLO3RyNa1JJJ9dZJNaOvhvdXmvczAO
e0Kxd4KNt4dW4ZJfCBe9QFgVPZ85rzah5Rtz4e6XV8XoCNzqK5jt68koLhWCLC3qCJlFP2rg7hO9
ta/ra6E6QyB6UGSPsnU8xSHz6vjmm1/1lskSQ/FkSDwp+lgGQxbhkqIqhQWba+29pA4PR48SD0CG
Xccm4rx/5GrRYpSkfk3jI905CaCAPxolU++avUGsNkWEfXyWAOTg0PoxAZp7T5prs3j2jhTIyvs+
yokBjEbtwOeSEa8da3usGnbaJ37CZZwVjB1B4ewjZ15ykp+MFhc3hmWVR1iwpmxfA0sFK3eV+iVX
mIxq+WAu7koG7lYPmz2athaBxAZf4bdoXXgUDi2oG2dtLiiZm5GoDOcuCLOdyTQf8jex3uTW3bHD
W6onhoU6T4sjjutjMKuyUNS1k2HZd426ABcd/ve+3GFnLDa3ljB1soxnX39HJxmuFdIS2p6p5dEb
V7fT4QS5mskoGiZwa/qYEYDPzpSwBXbHYKj9hYq8cQRv2sMxsu+QhYVLSIssxNVNQSdffbHgUc3d
WXk/glQdNnskWxqjufCiZI5/HNwCV/7s1YIdG0POPK442+1nJbYFApJVMWVzgSkjr/5z+KJJhBeG
lcQ25Ce0QyO3FXQYLXDTNfiMY9wbvxdkYMrJg+hnXDFWv1h1rYlv75/v5b/3nCnmM+fwyAp4kKJQ
pARaFYfoKX43qG3FuCQzpz/1Le07RHREgmN8kg9iJ0jIXNtnrz+xa9T066ErXlOV4HLXis+JRXtH
3cISed1PnjCVmOZGVwhLV1Jf63z5Tq+4HSh6i9aCAMUD7NfNtdvWwThWl+9sbbbL5cdwONMz2+ok
bfzrS9udntOPbPKmHsrLx+dZjXGHGJZNgzXgU1ben3zcPI2I7mpvH0mRc2rQ86+UxXiVabpE+X4=
`pragma protect end_protected
