// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lEIEGU5n+3lA6pKz939lxMjTlqjpEzei337mP9p6cmxZdpiLNQ60VKdlXaSZ361TVBCQBhugN2QU
bQq+B6yml1OwiMBG3wH2lPAvoBXBwhHbaU0BSNO6QFihILCHReHKxMPlELgRe5/Ot+PlbAAYk2G/
4eWmbu/GTGuJZD07wUzkLjp8eSjF5bV0HDT6JFmwkDS52MzbmYQPMOk+CG5D8Tq+k70Y9GSwD2/m
T5k6gl+ULE7ERC8POCdbFXMSgxArKG40NLDe1DYBYxPg48Y6AwrXRy6h+pQN0JbbtgIDTDRIHjAq
ZkFiGlYsjbhHPgVlUW+55jBv9JzwTqDAFp9H6g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
lPcDhVUIn25yNGh5HfBwcfvEAs2BfHx9NKMeJAeuAyYLCuMn7dBgEs5F1ED4y3oVSsDQn5I44n46
ejgUECjBf2xONfr6fdMRyrUUXhkIRtjekOLesfksAbFIN7N/12Yv5zp/Em6+M3D5RJNJ07mEduI6
QimnRg2oeCDC6dX30iyoUqkYud47T5sNng1nBMVnCDDlsvDBN4l5lSHpkE7uA1vtRR+anTo74UKv
rM7nHnsIo5KugEhN0AsbgqvmhH6Qrsh7Xdeu1KYHdzfE2teSl29frka9Ux5Dco4TUnAFP9pZO1Xg
8C+gYGaSMt1CguIT/qm9pLMmeYjBwYwkFOpVNcs7syh9QOYG5qp7GXE/6sfL8L3F95ASm6+WhHzN
uvPLOzOLpeZ3HL10gLU01vXtSHNbpn13wuTetN9CLj1bJpPg4D49Q+9Fs8pM9/dZ7J2IAL1QJ1YP
lGuTMQ3WYEl5eghVE3ZU/lShH4HYbE+DS8V4zTB4WbI8VDr2D0CS3uDjjZ5GGU8RhG8KOohtb73J
VmWmzCRi/cCup6tU5VtUBX9d60vlp+zUFHpsSVyjHpQSdTXGqLsY2dh9KFUYuC6PQdOEKnCOZ9lg
U2TNkeVvK2lZxGhh+FWG/IXin3WXvPpoHsjJxnvgJL7iEUItAnian6AqFHaooDy88Wl069V3JswI
3358ebyoj/VL4IoiJwxCPQFAWyeUccjszP6QhyJpo9DP2n7Di9g7711enFvfoUm36taMhNHc7i5N
lCStCfwMUlT8fP1XoNuZS2Au3+UqHu3cohf9FQEel3ydHJdbF5dnk1v6XoHcEtKHVFyHSAqdJoAi
wvlyC8g02+7kVwAEO+hmrw2F1cOnwXYgxFqUymWJNzq8YY3lzq5IgqWy4OfJSOLcvwpeTUi8nWoT
/hx5zpTSWCIrtb43RR+OXHN97Xj7E1zhQEOgxeZHkVFu3VdTwAOYl0bBXyNlpcBPuPedmdDb7Hr0
NQSFHnjVz817R1gzAKvkEDq6hlJ97YaovknshO52rh4GEwElcPeLRLzxmJZ45Kh4csfYmZOBCTwj
cZtEi7WS/YGdAQPfZfximkwIrhZ/yYsJSDC74lQApRYfM8EA2LCiF6SyptT0aFERYnsATKqagrA2
uRuNMb2DOcCyCFQJXt3mzEg0V0FxwvGMNNMXrjV4cgpUg3ESMPAZKaDgq3adbSpDkqN6p8EYN5Yb
l0JkRnBP1BvltmFOHUd3IzEo/aLC8ffTtpgXJOiV+yzI6BznA1xTSHoPH5Zgfwf/4R2fu7yf+/Pu
pU0JuQIZEuAbtp00xOPcXXrlzZlwQ5BDR9gvYeiECHiYGWNCliNjXUaY4f/xyNoTlATrio6Zj3Za
jStNXx+wJwrn8zsV9iAk+dRzsvgSWBo0NU28TK2mZpD1ZskpGzNjPMqnAi7RDIJt81+oICyzBaR0
SKUBPpaj4p+IxE35S8gmWe1i7Js2axH1q2UG68DILwCdzZJn1taIECmNifXgjMTX41kJbBR3srPL
2rdZmiA/PgL+v5w9r129OMfAlGynQ7immR7AeftSlc3jicShpCOoswA1m4QevE2x2SiO4HsvjOIK
YV5Oji5eWrkaCUU0MRR3EZ7vUGTsqGahfjBU0Mg5qGKuAJn+oQZsWli9I3whych4QxFsSFGZxez+
pb77ibv4cJO2UNamIMod6sDBR2XrYgOJCOtx9X5g/pjbp3IZ+ays6JDTPccusnucCvY1kDBifIkS
VZIR6VWeOmL/P2pZ866XPybn8iKwtqedYDaSs0rQDnfgNJnPAIq2YaIMsR/QqQ14QqiEj7J7k+5p
HqAZcLbBOQZNXt9hc7uWHK334Q4YOo7jcRpDaDiF8DhfqVkySL5bVyl5baRwHQFkLqtUz6QzhBJe
8wo7wbkIm06tJVFR4L5j/qh0Co+Ma5ynAqxxJ084vqVBLItMBUjS6Jk+OwVD2WHkIpz9KzKpExS5
ZJL2WomtDTHqCzMUkN0Byw3JHkbh0418QoBfugiyGosfpxWYWNBm2WJZJ2ZXJqe4p980NqHKKH9k
O+lUqhKZ7OkNtOydWK2wjuHhenM9Ia0mPA/8oL973ZzYBfPnENcdMWxpZxCTjG7Y6HplTeuVzv3X
aweJLtXdwq35p++9AvIQqQ65ffi1Cz/+s5NCq6OLMa1/UdRShcBuqUeHr7Y94iKY2PwiPVMXbyvP
VaUxJrdMA1twkTSKZ6+yrUdY+W+QInIQ6beLgNQVld7bA4nSeMUUS9DNZxVwQ5RoKOSJXE7DPpLW
LWYyZ38qRJQ9FyX2u5bKIX+JyUlX9YFJTs31vlM/0pYsTm+BUSBZ2aAHOPGXtTxVGxWvUI73vWM4
XOMubPyEr5pn0rLTdybOb//2rTEcBJMPl35VUCYevmTQh/2T4iUIXJqRY7zijVHXRNIgGxivqyZA
lvpStyussz2DviCy418OrIIUzEjTmiWifchhVcO/gnF6wEf7OsGs2f1U21PBruWcQAjLb2+F2h/w
oU/y6QBwCbaaf6I+cmUUoLi82893lqRDq6qctbG42QqnAv9uR7lAJHuLEoJTXX1Osx5JVt41/sI8
wEHpIcHhM+jDMNPxKAyeOw2qvUd0qEoJFjEvIoRKB+WsHHQ5UVqV+1915LejkUCBk5ABXXwDUepu
6aF6mbldZYOWCG78peP7D7uMPxDW93kZEu+OUhgfkecdKX4P2J0Lx2GLy39zxe3Bhi5+Ts9jk0I0
DmcFkyEadeMDOSJXSKdNoMUobRcP3xxlowl5vUhiWiJ/u4wiv0cNFhlqKLZxOXoIKgv9BKYmy1FU
JvfhShSAGENX1pJGlPlojduy8SGyR1q2Rx9FUeoKfYRi+0WnKEE3SdV4GqGj8piGbxqG6TYbgCfu
8cZM5azcFHlcoaIDfMJeKzMQfbVsAQpJdZpKFGZV+CLtOkj0CDJ+okbeIuZa9CHglcNinJyUfiLF
1qoF3L2nlIGYprYJ/qoTGBLaC3vIYuiMb4bV68AqDeBjnEwg8IYgXJXtB1s5qS+M5uwNSFxEuo2I
UjNckqoiDr1Z5RXQAz2VpPqBTz15+f9PykIBuAHjyvUbOIx0wwxrzhFU8eQCIMQ22vKGsijKI0h7
opAtb+au3pd/2bnnlfNywscuslukbwScBCCX7Ml2PEWEKQ+mIYfkF2wf11TgmA/n4WGj1r1yxCuQ
ff596423Rt44MbV2xzoC+1bc0PNY/yJr1NWxti9XUCQMRg+YO/VdF7QkxdwUuxQQeD8GSRbuFPMv
FIbgn+HGuD9bhFsoPpUWXnJCfa1y0O7GyPvC0UB5RfntACOJTBB/V/D/a2xWw9aQY2Gm5JvKhwjN
Ce/A4OROMAOou7roL4OGD9a9FKi7jc37PFXsiEz8Of1tJoFVxTOXSyw3fn+VMlx9qrxDKRxHVbCt
ligKpiLagE3dLOPH2iDP/v7rHQ77aPj2msQZRh+X5F2d+P6zkRt/XO0dZdfJ8JOP+wZKiHBybzRk
YXEMZgKZl5CXY8oiqldIJQuMDEk79pQrJkn2c+JererjAm2pSjmNyyWY2FOB2mZN+lMimBaCElwW
P+6/DCnKsul5wGn/UOcAf6urAD86QIVsyT/t+lr0O7td7UERe5+N5o7E4sV9pT/kn0/03sE49Hn7
auMQ9MvIsMwJvNqRtiFyFUzJM8OPUy7mUUI7Ai5XTbp4zHtZwTOFhSsj5JENo5QoEiUweBbIIzLj
nap/7ViN3AjHie3fdFRw0DgUClvBgFhwkA4YpWch8D8nf/+w7QdEGRh50MSi1Cxg8iezfAQu6aql
TnW19LyA7urpJblxD9FNZLd/jpxq2tfm/Q0Q4rSWvu84gKJADXskrLxe64uNftCDqK/fEzxIsZ3d
TI6kfdYlVnDqW4DPepA/n84EmQRS6qkSAsuwmkwTEcSXJZlTAbrkUI0gbJ+CQ5Gqsb0xM6Vg/yVl
aAGxffYEgVIBUSjGYxZNCcOSRYt++fz0+uMhT+KvQtjn15s0jV1Wolx7wZrw5T+m1VSXIBKkSag0
XUJ6ycdP9J6/nWX2hq3dUJSuP6kKjko0OlUE/v/ovacPU3eQ9ChTa5W+hs5YipBTuY448PaLVdW9
gmMvLKLivIVoRY1tknMWHLn9pQQmOGTg97hUGjtNeybt6FNofdtjqMuA9E6oHnDp+a0aJjcLk8Zw
42xBGguXiNWkCjc2GE+T6byUXnt8s9FZWY1glnP9KVi/PTNSDjkuK4z3mTZJhkJlHTZvspP9NeAX
BlK5EiJLtz7vzh0Tn++tAzvGd/JU1YOsdM3ZwzdXbmLa2TpX6ejDulZoEWOygC++kQGzFPyIvF8Y
dKSw6sPh2+8ijIz5YNUJjk1jDvuMcZi8am4w6GB6oBvz/PViEPEby0emGIUwsHa+jGFeB0bxqD4x
v1n7Jk7EjNVHjpqfMs+FrvPVZkSfJU+l85Fhtpz/UxhQ/y2Lw0KXzqWf5BpwQtoAxLRhUfFD16di
VXL/daZSM0YmqOeUow5HqV94WublECezl5c4w7xstwmLi/QBhZoL9H/J612C0YzYYQHvj04oBPu7
Xbw08eIgTBn0VDiUG6xfEfiFcvRhx+DEy8+5td7J4Mdku0Cb5Cnws6X3GvUFlQ1p0CPrgkrzY1P6
SqRqwWK1dQPZcVQXcWoQqT+zoHPbXq0gP0fOMOQGDm8MZWgkqcSM0pJ17B4kBuBuA6MM7nfzEkOp
pc6iZBOYPJa/ELptmJFMQRgJukVO4Nr0unv2J5KsX2KXGIALt/Wlvk7OxT/R2c8l5IDG4AmIMnP7
cD+Tck10/oPj124dc2xKbewIKnJDZlsuM5CmzwRe2gMwGbtyf3QJLF4iwgXpmKKK7TFkOpaOX6Di
8HEBMAGgPRpSYo4m/sr901QmjjHeYzj07cViCITjKn1ns5XkHr1fN/Z6wQjuKoDXygeEmWjiPkrb
hMadNQ6sKXQRWsB3XjEj3v5Ivlv7leikD7CfW98PPb70Dl2hvrkvtiH6T/B6de7iPJh/NUEJX6K9
L9QiGug4mxw1POfK/3A3qT9oVbnQDkVjy0kxx5BDgU8jUD54Pf4a6gUikvTwZ7J/8KSkgOBOpW/+
8kQhpbNUiT6+QFyyHPEvqsfXwrWr15W3bJcemnG4gojVAW2clm5shHKruPrfjbk4vw9w17qnWVzm
rbE9a+RfBCEQtcZgao5vfKpHx6DrxD9llOIJpLF5T7jVeT2bQkjPsVHA/UdzwcvqzgMxnbP8xYeI
v2JTy6LLcgSwMonIgfTRHN1x+oQnFoTS4UxdUtpK34FE/xAyij+89ucgqfSjvvkhYazR2xx6OZCg
lVwSQiQd9vB4vxOI7lfAur1Kv1aqeFTUkbDooh4ZVk5G4cfc6rOwFkjVmDj/kFkOe8NMswl6DBKq
h0i1nFHAg366l4ViuC3lDrAXxAFX9wt6sj7fe608R035xMQTLHO6RUlwRaq5hqT5ukmHuqKhi8xo
Xp+M4LggFnnLoNwpJbhcyu3tjh3xquOCsPj5iQoJSinbsxz9+l0svdVxJyYSVeHSMa5GOifvOUCe
gcE9olNnTfLnXUlXddDdjOfhYMHBPFR8bcafhLNMuscXeU6M4kRmL/pxaMLjAx98zTbWHKo+tTvx
aiNowvPW9xfNG+nX9shwjYr/HPtNl5TpFsut2FaWCDOnrqx4EbTA1u06hk5/g4BJFJMyroPIO+iY
SoClrTWkTx8BpOwqH/cKn6CG19yvjs+tWMZpqX0Qw7LPAtc4eTp454uifnbRG1WZsxLsbtc3vdqy
RMCazPRhCaVTa8qSPf+DIPP4u1MYUESVXa+HZBlh9FZua40eMLheIHXdAiImafxwQ4PNBmB8Z46Y
uYuYyUjLo2n5G0oPLQzyHffdN2zFwZcZCFmDUbGtj/3YDO1j0KCq5yZT8u597irZxgJ3prbbK6Km
XyjPcMCNMFG51a6EtiPoD7pDIdZLUlrD+8h1I9u96RX3v8zEt3seG0DPGSWT33Xm8/qlPoiNp9as
RRk31gZCNChg3WtXxPLE0YQPnoBILEgjzmICEcD/xf6tg8SUKbFGwEKEdIbsTZou/npYQlmi5uwh
E+tSyeXSiSxdSMhFsVfM2sYHszVxTOVgev5DYvg9dzrt1Z9xwmx0ov0dp0UicczKdCs6CqsvYmTv
3LRskOEPHfNxaQEGr1b9lIXkRfj+jxcY5cF2u1pqDykEGleJaevX2dQG3DjDsnItIK+byOOWYt4P
mhdh2t/E+yj1ayVW9u+U4zOEtGG6GuUEz8rvxYU2zhN0TnqxHQpmYQn0MNWJV7/MRerbXgSCbFF8
6sR6oSb/bIZ+tAd54TgqZfWtSDagZi2yt86ORyrR2yLUU66R7YFTYQx3YaVSbGcORdCiGJEc2smE
2Zf4ESAJds31C+ccDNa0K8RBNP58NbSEgYULhq7rg2Hg8z72A6VBTESCjpHpeNRyI7JbOWhWwl/N
LBgK9wOLA1LQiYek6tmHMq5bO+yoAVLI0YZEAhtRWJkCZwPDkUQpMrhYUbapthjjInFI1bJMw1yR
ewjBkQn3qA+FZFWaTurr6Bmd0jUtE1r7I+rVzROIpH8dhvjGp7x6hbb/BImISOVGdmWMOEduo91D
EeYKRDDDeZ0cwtxsxa7oz3CD2phw0ZZ8Abi82Rb2Pdhe+wyiw4vzfbGuiHPbcg4yijd6vigbnA5B
pZ8oSXeXlmp8JwVBIt5kFCatcmtUyIJSlNw9Y+0TuwnPpzARu1gP2WoxQUwXFe3VsBf57rrpgfTx
5E4qjf9ThgSt5tLMF2tQTL3Zb7LKhHQk0GgVScSRXuicuDQVGw3Uit9tKPvHIgxrW2lcLK/+3TQl
BWzL9w6nisHkSeFs7mfd4Y5c51ZG+viTxwf7DsrNZN6ieaqmjx28uHsKFuloeGhtJc31CtW6Z/er
Jx4jGX6trhoiXqbF8vBXLUk94QFwpQIotN89rYlvxdAwDEBMPTj6WXrggSCHS/Kbf3sJ3OgfSu9P
pEUliAIf8nqRkZ+klbBS/qMtMrdEKtHe1aOf35hwSR3ha3iSfypKA4haOleIDV46IbUhQ7ije7mI
v347536xJCHDvtuxedh1SFAeQcoQvGouLqw2JszwIPp2dP1AEuDPdXDskNSxh1w0JOvNYZEMlHBK
CokbPE4yQnQis0ps3WnsOX86clE4J1Qk3kTDR/xXuU9ZVoyGu9YzTRYkdd1Opdm/+KbP06/eyBTc
XUA8+cQ3SlFcO2MLDSvy7cyBIaktHXoMPaInDUYojP+N32Oka6l6tlYvjQU0PfzCvAYRBFeVN/7t
eXcyb1waGbbG83OEYdX/BvmjyAU4suR7cKL6BlR7bvHSgauFFJn3fo3SvaTBRd4hYa54XXy/mClk
p2rsWEdoMt1DqIld+fnIDndLNeFjJ4h5VWYAxMQzPvTaZhaZMP+VkzZpbHIPkEpSm+fEEN3a7J+q
c4E9a3a5rcICu0NzZ+AM4FoEoKg43IbwX/i9qY59M5F2pFGAkYO8Qob0lh+EKWdMiL+JgcQf0wON
dIrv93QJ7rrG5FSMFyPGBwkraqZEI5WWkpvMtoGol8H0Qo7T0f7K4TIDgrI2r0wongnnzYIoQx/w
QbbhKdO9NhrfhogZU5MuWQ66oZH2ZkFnfHF9e7lmaHdKahvrzmC6lCe9mg4/M/aDfvQTJBcvU/1g
IA8Pufog7yvLOAlMgNfZl+Gij2c101v8rqHjxVwGWXxSD3vsn9J9kIg3wIxuhGBKmRe8vN0+SolH
AV2a6Nw6v7f0pMQAxPnK8/yeMDyjWg+k6JqqMsOGOKPHN7Z50r0zAvXZiTzqgNQyo5GNrH+CexT5
0Cgxit1Aht5GpMdw42SYK2ytc6gqS+AAnJEMt12vQlZpRa6FnYWgvfdGMPDIUXujzxJVMcN7GSy1
tJZWRh2fylXWXwKZC/6pt1D7uHl4dhD2yV69qo+kgeqhDELdRdt1IcOOPdVmPQOCHGFpKdZBL9rK
BgKQYhtSEH66Rck1QYyH6Lld2/rKBrMdFm0DcmTb7kKe1e8oopLOSHUgu3ua+fLkFcQYHeQGIBlB
vT0dl/zVTwS4sl6b4e+cYbaFFoqIG87A17OkNOlhoJXygBhJWSVzHhemh5LplYUbjc3noyZFqbSO
fzEI0hABaDr1ALlnphB8rLOWR6ce6UFGRXtIRIOX0J7qM0S5YrCwR9bashDakJAw3cIgPKtQhXGQ
aVF7eZmnSvigwN4ML6BkFXDbYsVJMJG42y12B5KRt6UMACU/Ib+t2/+CZhiQXaJLNxsJtrAUuFmm
A8R6oZrr9Y2gqG0LmiL9P/+zLbXIopSpR69F4H19TTimF7NM8YR5BWTXKoaeVR13Kap6fTVe1m6L
FX8iFgx8g14EL4woaIYYZaVtgtJyVrV8dAhONlAYaC/A7GImVuQhLyAOiN6zPtDWOypZakcYnph2
dIXiVkKz7eEd+T1Pqyq0FCwGV4i15dDtm5Yn1A7H5dBsR8kDp9Rkt3mZgrT5yKuC8qeKaLx8eW1f
2W5IWZIS2A4k46n1MvgZMSQ8sFKfhvN+f5A7lPiImJZFKldnYFtvAKZ3ndPVN8RL3Pex4sX2+wsE
9iTuEEHPnTKpOb+9kFFc8a/GlAwgZL5+PfEIZiU1ABdmW40ARpD332pfsZK3CYWl+RZqH+QFQbE1
sQejHmLOPe4hf9EvFs8I8+e5XrqMZAQl7OcJkz7dV9CR4M33eaEw0MhvDkL6EQ0WmKPDipEZvUmy
70258N/s05dEyzMJNuF8svFBNh9CtNOF3Jnm4RtvDaga7y529vt20JqWhlKAkfo6IhCgb2xVCvbN
dqwFxSeVVmp6JLALgP6vvY4Y6O36uYDg12mFaqIg20Mfw1KcDQVu61kuNeinChcJdpNU800Y1D1l
WCxn0vXgTpXJuxx+aC2n24E93RWv/xM4rFdETet+SzpmAaa4aoui4V+XCS78IUQO1aOCG6iq/5jf
w/HE0PMK9KfwxUxfFKAGiXMTNjr/sdEYIB8HvDUDN8KCiMLWgCKTvqQW7CGwxNeAMH1pCw2UDssM
7I9/N8nJQMSbHCpZhJ8KCAxTwGVp4Z7i8mPneVT24Tx0Ar+6xvZxBzy5fI8/TNBQgVli+TckxcBZ
kC23Bhv1y2B5v4QHgzt8rSNOC1IIHQXE/lDujJaGtzWffGSqtMtsmnn5Y9+YK/jFbzSjDX5CkKES
k6GKZ3qQj40Bx5nspHDV174nF9Y1bMosxEA+6xyZXiZatIu+mh6zD1tD8Z4mKyD5+P/MO8T7ipKW
7vswmNcdsA4DUA/ph+SyPEhgGpY49YnoJ2RvdCVDi8b+8zUciQer784UjQvDI/b5f2w6DaVdtRAY
GzJfznj5yh6TBuqPjSlR1N2hEF1TkSctl86Dm61nnNjryaT3e38VLbn0p2BLz+y5U1QxvtejiRdV
FNfbWWTffxP7+1wDb8pdO3CzHdxP5uPVuXi+I7AsRnwx40i4XxMqGCZ5Jb0MI/ILexAU/5rUCkOb
fS5gnXEDFLDoVgV7aam7aJTZsp23BZs3fx5crU6gxl7NemzOzjRmVnEKftdG+x5ALTiUlND+OH7O
p3nA9JTMzykqwn1xf3gowQza2iu7ySQPR6RYX8ZMQ4DlelkjWDCovjf9V9pQgDd+BQ+p2zrvXp1S
ossHwWlkYwj8vp5wy7/ceCykzWZnmFwg7U00m1RiiWWrk4hIQjO4jZyFjl6nvevkSX0L1EmcFbzg
NoaOxPGIxYIYA9vbHhL1JkgaQAgrFbBCbnIrp4503dsY2f/PoMHFmUVgKQsJnC2ksbKRqliY+8mx
B0Y8nY83dVD1gWs4KYkzcJZmHmspaTRelNbhIbhvYQ8UArsVQrfYF+Axc8Q+q53KY0zoYt3KX3r9
2tGeajKLh7vaCK+qNV3Ob/j68YxknwxXVvaz2TaiYp8dyRgK7qzkUiSw8bW8QVXRlMwYRbEwv0Pw
wj2IJzw9yjukR8Qrd/bECVMMYHhonqZX4oy3DNfrRD3dY/CNGGjAYZ/FHT4qCbPP3x3zst4Y5GQb
ITyFJSjECn+0myg7rtxttQQPoaG0YC1TWcCUETneu7TpRHOXggDLIGZk4TwwFT3oSJihvwQ0meRk
PtAET4xlcrG745zQ+o+Tfku9hXaadBySV7kUpIgqf+m7klRjfOJh3B48W767HuQvpbPnaq4dg4Rz
g/r4hzuN1utC453rofA/V7ep1u87Dhh1dibHXUMYTDbK1XFvBgMQ7m7d468Vn39AE6FjwV1vPmC4
TjZwnwU5uVrH+m2lgcKBvc/mNfVW1m+vA7dwOfJTCT3d7vRda5tLXk96HHe6i83DkIcPAVw3gOpo
4wedeqwq1kczwRIc1+opc5IyroBuw5bBjYSJ7QE1go8ACt+bnI0R7r5A7oMWajJS798j3nsazIFu
bIvzAnukMWDKeRAengLTs3YODFiTSdRaMlcSx5SqU1CNylOSoYv9tpd0Ib0RVwJNWonAsia9wkIf
SFfY9LacF0ptaH0ZppNsSmSr7aGZZPi6liUBt9jDsqAPp7bPX7VQcbBDyAax95QG0CvN2Bt8tA9Y
4oOuJcgrLoGmi9+t9VLKCxRcZHyHhbIvVHKHwoBsqiYO+5e7HYw9rqnBoIvG+ip5FkUFj+uSYehs
XQwm4AkEtClwYYp7eDC4PXY4wtwN8zrh49ujCo6WGs798YbsClyZrwOITa90qEapGk4ACnDb5byw
oboWqTfRtc0Xwuo8Ws84VQUlC+tW2JshqUVvZMMCh5SWkqboBzmOvX0c/uOFK4XbZnqszPond6kT
NrS17b/CO0/0T8LFu8ciPWEdQhD+8r1I1zDnMX4Cl/zwkuIJT14/joxPTEeKGMsqgY5sommq8o9f
ppE9NHTIzRRGjuh7Zyap1GIyGA2GWNaLDVyrz4uMoJ44XPljJnd7aR4VvtOr5sHIR+NmDx8D/3bk
KpRyVxvQj7vJjcm2lcBXhtmg2Ij0MUSnQQ6y9IdsiSd3l1n38ogBkkmbWySvmmtsMNqxqMNnh+se
ViqjJqXRm9vhbG9inXZTr/TC6JhsG5jZyoiVLaN8JIFteo14vPRJPzfzo81AEEGk1PgqSYais3B2
SFTMtMqH/qHxC324QlvM2ywlpBemQG3l6SAeFETcaTLEf4Yx+Wd8rtnrFEOMegjIPRt5sR12fa9x
MXuiJg5RFkK6zV00P3qiHjB3q/egHFWlbZH8RBFlzgszRc6YjjxHJDcTmEBKphCBX+VwaMK7Lh8v
HO3wLEEPRSC8A2LOe77/Ixng197QC5cDCZIUrhwtP+rm65kg6VU2K6yZXh8+/eQH6PpaW8o17zDv
sioWb7iPxVI9kS1L7JMiY4GmA9mKYUUjiw2csbJ4KMocbtJWXHaD29KRPC1NPMpzOHog7CSyQmuq
JEElJqXVYdFh0eSqyNRejyA6GLlAdqAj3150jMYas580K31FYjEp5rnLkwuK7hcCw8eKE/fR9SAp
ZKFUkALqav0OZWpH1h+MG2+T7RMc7Q0LzTjvBlUO03z8tnq7VpyOu0X1EKNjRYpKUbykJ3aENHn1
H82li7liCHC8jNCNmZGO+9n44kqQU5ZKlAH9UKMRE/DdtZna5XerrJi1ulzYaZcZq0pk7J1qDdy8
iN2bc6OB9Nz95OMUus92xvisCKLTKjbA0JnvIszle4PeqC47OyOPia5/FN0AFQ3bLVD8S6qB9h9E
g1FTWartkXhnwh576tj1qtE4CuONrV6/cZWWmUwgxLJlhubfBCtIuFxk6iJpZQfo30i1dcQeeenM
9yIi8CAZ8Tt9lf9sZUkWxDOUc9VaBW8MMzEa4QcjwjbJWaAYoPuoFX8dFj0aXZ/xTmZqWKP2TMjX
qfOpXPT7DK1Ro5TA9bWsX+1h2Qck1Bjy8skFzfBhwrSj04kiwAXqMdAKYPtE6OTFZP3wWHwbJxHc
2G7PcgXmobR66dhu5TQYo+FeYac5Wtd7ct9j5e0njklPgpmhXKilmXGO7b8mCSdyoqI59TX1EaAY
x+jJQa/5H3xZQzmC88tsB+VkUhRJ+/gX0djrt4aQHEo2nWZGQPhK6WrrZ0pTYfQQHKbmz2IqkhLP
fp4asVvCbmhPWqyBQca8+oLbvNxAGQxlvM9hvcnj8VTrnda7Pc8WPO6yQtEiTOavm5WSSUCkcSJ4
F4WMF3NhwQ55mc3lHzD49PTerA/afWD9gZcK+HNHzJIpD8JKSuJxMhvn9Xyppyi+lbuQyhbB3vNg
OkmWxMuroTWcYK/HFCha3e47FDSIDGoBqmwbRp2QEUA+QZmx4pS6uoggLn3/SrYKxmrRe4+/G6zE
Mb0/l9FnomEGf9bU7noQpI6Ll4WyU6ib5OlRoDe5WBGq/9CfhQcyx+1/FHOQMDE5gyIbtZ82EXBf
1S4nnN62IZGSfAP6kofj7UHFHem8PgWewe1chzTuWrsTMlF4nwKjHYrRYX8V7xH30v2f1IcOu5BA
7ku4r42T0Ems4LdW68nGpykWYXjTS2fEKiCq6tZorta2+iyxL552tqQjb/eTaqqIuvy3egnDFu8F
h7noQtxIASMO9eUbwkW11h8euiD1Gqtn6UFbsJMta/Hic1cjDvphr6+62DwUpoxUyC4D+FuVwz4y
Xv4LGocGG34qOC/qQRRyo+l7cxW5DkXaJGn6AZb/qnTiXWYymvt+J+QTd2a7Fx4x90PQHKoMV3AP
13UaSiKnIbFmJ/kI1PGBFgQAfAQzVN0SJ+7rCImnPGS027qwMtbjrXpLaeCYaE2XrTj1CyVhFOCX
oXEEXguHO0wlYAr0HHi1gsPsTKrAMEBRfwxeYtCt2OErihBhedTpK3N+aMNbLIitb5ZnM0Q6QF20
JohwN4WaQKsFlPjOiKhav7oCQsLEcvPD+sJwr0b0FluquTq4qyaZN0S+S5w6nKkNRrAw7zY45x3M
AvEKTnr5entyUz7Kbzo5gT7r1vLzdbucdd4wxVE34RhicWgyZIgtvykPuLDvudsOECdDVyON6FL9
G6aadDqxjBXaobvXvSQRAwJZ9vAf+7AYrNAcGK+q/RPu8VzL9LPIHt+Z/UI4zRGdvh9IoA1fjGs0
CQVTBMTHvts1WlKJwZw91axhF/vWLpoZD0DHm4xbY0Q/R9VKaDm4X+TdpsqX2VdacOk48Ab4/VuD
98cWvHcbq2hyHr59edst6gzcT6p2LWl4RtV+kWOuivrOp7hmj5npgztjJwP5zVwU/WFZxsx0JHjf
z6qT8285494NwSt33Hrt9+1ZTebt0bnWRlN7rTpEls2Ef8Jbpzozl2nSJVZMNIEkC0vh1j42ty2Y
WXiJXQ7W3klV/e/lJM1T26TeFLgDYpPSyGG8n1AQVjT+xC/zQOxlEzT+Yb4o1JUx4HbEjnXTD3Wm
uHjPVjyl0rqArGhfjiX6Gi5KbldwaIjW+XZrhRuzEtN745UVJxK9XsiTBLhFYC0BBQngh+SoQcEe
bv5Imr+e/S1uTtcEINUuw1fyaA1gAPkCb5ZUi4CRix6CUZq1cSC0qq8zaOzAqmkDcRX44ykO/Prr
UQQYQqFqeKtXEQlq/jKNoC3u0gUmbTkWyDbyBR/fO9hT3uaFfk5jBUMCVnrBXwdUqfrEzQ00SUm7
ehzIXiakZ0v78xrVq5MyhBHeOLz4mWCsG59q1Hcsv3sc5oq2FAjdMKEuiud8I6aK3gDh2iRbmd8h
SjVJxiirOFYz8bNSMt06L4c71IrURwC1QmAC1AL9n/ZKu8/QonDbKLHntqr8Jjd9znvnfcVfbi0c
O2shSblHoyDp/GcB2OWbWrEU7lCjGzCfap0/FnP1sECbgySo7E0wwpnVFfB7gshY36QTjbYqlJxI
1QGlAfueauN2cYujL+F7ppXO1/3rHrjGkfklpvYLeeA9HIyNGvrPP+1H8wzgM+QOhATwskHHG+za
bB7flGzpV2uyrL3m7rftWmWoLaBmeB0mDhU7jJ/n2JlFSVTbyHUokjE4z7oxNSSQlbVu1OMD8bKh
9+BkPpRSh9z/MU5yxSYDW4HWVJ4MqmobFn+gcdqf0TEzThlH7+kqWEDrWAROb79ccrjAatjqUgcL
ShXUoC07Mm20GU/4EHP+f9u/uGz0cF9q87WA908hn+yIP5oFPpRphY0YTEq2EDpRC28sBU1C4X/r
hlFiQaCazaJPxVMHp2Lp9bvstp+jiQqEIpjEbB24IOYEdSjaS7AgsHOkQnfk3cmrswhXhMfobCZw
fkulxrNhtjfn2r5dhR+4cZV1LtqbroA280FiFwQHGGwVh1OoUftM7BBJ8g2g9pktD/HEf4H6skq6
pKz/5fONIFJaIq4pMZ8oxQKVN6GhlSI2LYlJvSfarBiebFSO4WA6KV0hT4Q287Wf4Ima9r2S9IQD
xBBFmwo6RMNCWQvZU1//oEOS/h5D1BmMDcpNjD9YbKUcOFpBfrfx+sA1sfGPiUMwMVLNTrNrRpgl
1uSg37/9PxANfzd2zYtQDnEw6ihJ6IID1p/lJYm2lA8JtzkVJ5uSA3j+lVlKAwqfZ9W0o8RmpXYO
9iD4T+B6tvYJZjvlrT6j4cvR+JSI7DrhAC4kRoUgArRj2nhpo8lgsU4Bk7WCYTTyUvgo33ehZmyJ
cfJFCe+DcyuDwO1MPh6bTfxQbswpD3Ho6JNbzSatMX8kkvnRmDR0QO0ybtjABrutxNJio1p+J5pV
HfknbvF1FtJeaLAaODV0xqQo7XyPEtRwcVrk1lvzZk55OrDKsIrItXDG4KNMFFuWGQZmI7BEKvFg
in3CDKCxaeK9ZaCufkSXvYpFjD83qP+DpUfoyy5VLUJ0F+5kBnG9BCTWnNiQkLUs6xgeRaqBjVx1
sXz9O8n4e6lom+fqDPUQhM4X0NRBRtCrVMI8MatXfoCaBmMZwmCo+lGQs8tCqwVH+aQEeBnZsowx
S22E41WZjp5/jGXVACVHtlWn4zwA2v9nvVzzj2xm64TnNj7af97kT8tFFsqI5xJJczkxoV6L7+Mt
z0ixUKWLK3L1mcsbZJmiCZide0SXKnE0gK3ozBQgtgAqJtRYfGwttvQwECfVO972JeZLbM+E3liA
EestyTj85r8YoEF2BX3rn88Vu8lr/NlnrsPJtkc+6wSidkN7ef9mh0d4tFR0nClEC3YVQNCO/q5k
BzbhgGq29Fu33JyYYD3gH0Xlr0ZiKlt2GmZjk5JdrQhtMecDTHA2gdsyyiVUpca5OSEYFcXUBqg3
Cu094H0cZ9VaKdoHbZOfcBxAZxoJLSXBTSvQyzgxnENaiZAUWKjTkUFdAHEKcTsA7twgnFWuVj41
HdoNBArEvybLDAspQcw8m/ObxoaFwh2AnKeyTlGFeGgcAam76PKDfR4wW+tLUQrXlc9GtnvPm1cS
Aoy1nevycgI4TXvkdTcnDtv3D+YmL4Emn1oZ01dgGu7W+C8WN+ESsJCrZBsOdyfLDSxXDZPXFov9
TCH3mRhZrWOPrZUFLo1ZWWUK81qMWETaHW5ai4spaYCXM9pahG9RhZNEFds/S6onlPcFVKxr+RBS
ZOrWyMHQyMBAB/3sKRo/KyzH1tnfMuZx7gj277k0ztZDuNKZmonNiowwwlhq/TZgDrsC0vrROOyH
X+F7h9G4O1SY4UOp0FulOWZMWhf1YerQJeVspsR/fIY/W9AK3uV1OWGrjdqXSzYMlFTRFkTFNykq
i9gjfta5EBLYCyHyaoxe5+E+cvfduE7GaTl3pT0PKPoibzWmW+IKfYYMl4vWXVMz/AQ+90LVoAMn
07nK0IApRHoEN2Py0HW3HCbd1EJIPBn5UnHe8HzIgYr/x4LA1914j3nRTduKQHcMevpvUgUPAsKS
V8rclXCxCs7H5NJuT7zkAjWCOfdtA3p2nmy5dQXyiBAT/fG/ZeTS4DVkaX0MTodQEdgG9tDHfjWV
EbiVvxHnoKH1jetdtoi/z1/9IBsiUmpsSVCux7Si3peYKBNNYm/960IgQnQ9HMvUCPpRibHA9y4h
MPwRM6eAY+3sEad041x85G7dGQM8RGk6+kGHn+ZEpivHwExLYUDXyk02mdXsduIzYatL5Rs8Pci5
fymT7YXJFZcgyVp2kZfxG/BFsfvW5kFiJ8MeRxdhZu1fmxQZpHMUoeS2OTYMnARFtsUayXv/v10S
ReJRJ3Yo7FQtjQksljO6xYk9dJeaXrhpXmywscfta1hTpo7R5qZHngrfL6dqP8whHWqw0VDtDYrz
dNyfwRCWa6g/BicNJVfaWef99xukXnZNFX2FQ34Jja4Mz2bdF8dXrEbB9syQFhrotAtEaxXSywZE
nVI6U6lpznN7lVAJ8Wqvq9rdVVPICLTx8jM/KUXKdGywwEdjnPjEw7tIrUXY8Aj0cIegN2uuUlqf
D9KyFyqJh9knRjT3ajGtGqEqRqMAHokEapN7K/UjKKSkmZkDrBubyMD4a76Pz9NLYgOXwoaAnokP
26IhaVfgnLfbfIAoAUr5KVIzfKONSlyWEj9rUodfGBo04gtZQP7IdxMzx1baMpJdDH7niZP4PbJe
vpZu0umsITYupES+uLgRkvMaM/Xr2/t9xcch2Mu3kc2aB7ITqhUUofPe2fYK4OHIhVrgc+/DPUti
DQzb9JP8iIq8uDZzvNE3i0PP4tYnxAojv80I2S5OKqhc0Cg8O0hZuQQBK/7SJfYvSABNR6wNkEIq
mnpBcZ2cmqQnUAknyAkw6Y4fqNPLQP8zCEtQT54jgTxVFahux2rXGKlwudJgTuLOg9ANyS4/ly4M
sGgjMLUEz6dNHMJFuhpFoAMKnmWoyX7zw/8ComI0Q9l79inId3EtV4PlJQ1fAgX9TW5mNW/4Hz5n
0lN0xztAaHHqvEZ7ueayaQH4yQV5I+bq+OwoaD3nb669ixpYsEg+8Q8J4Iv0HUTtK81ouYKkv3Fu
DEzqnm8kpn/L7O0YAqGasPLLNpQgTEUP8/e/wc5WOFWSW2Lvg4Hsk1VdYcJ7FN1I7KAp7sOOXHDs
EmeIn7YSJrhovG3Zhddsj1nurKAkesJIwPsl6b9t0feUOkud0fzKHiIlIYRFx8/2uwNhiZ0AogFi
ujnFhIY0iNaeSRZSrEDPEifY9iLQBelaHsD1tKEcM/o+rI09K1tjtU5jrSfeJmCu9adjhxBq1BLY
Ypx9qI0gVOrNww4P5aHY+z3oaDqm28GRZYRU6kxRwYxfhQ7DTEkPeHQvA0jwP5cWs5wFP4uLGrIU
F3KSpmnfqvbn5MH6NO0sCFhulxAiqwXRl0AH5wl1pOTpSVmh41rT4d67r75zarqNP5Qf3LLL/yq/
ZLuTQ5K9J0U8TMr/hvlfqFL7ZTLFxVhCGS/1rjsAqGnwRd1G379AfxMA7Y1mZvtkTwnzrh1KXmqx
XSdwpBuZSVeBn5B+4dvE2Begw6LQJLy0ZgS3rxZmVDGxJTvUoTgGN5GbWhOqi4r1vGK1f5nkePlq
/lV3+3gC0cq4Lz1iIGhPcdd92NVw5+bm8tUUtAz6WL21qd+W601vDaknpVAGrnB0twfZ11bZa1qF
TEkGjlufEpFCfK9agmbB0Pov/7A60XOStGDoGIt5abLHJk1USpEtSi4e4Thu4JaRI+4pOO2016XP
67fO4tgjJ+sSQA/gG4RdUCpGn7PAEKuSF/E5AeGIizPnDTyzJhFbDzcRWA7yv3akS5I79v4oYEoH
oFYXunEd+7CTAsrVNdqR7inwTKg+m05x/zbJlsRPd2EfBicyw+3OE/kQEtY7o7RMIZDY75yRRxhZ
VbAhpe42/SbZQIAkSb9V4lIqlvfnkFvkzNSaSWLfVwBmjyX9zzA5SlTmOs+/oiMVotz/gh26hgQo
8oahdPIJV/Wzh08gAlPRtJdTi6s1smrFDveEVeo3WSCTADHIovfjXW2oav1VlNtKDw4JeI07WUYw
zDvDjoy+/oc8yP1KcoFEjofec1M6jrU/k7dsQa1j+R5j1urYyvCeTZ+jsMt6zsDo3nGTXyjsIsCn
has31HuloNDmJhSPjsN7bfnfnhayiM/3SZ1Ph9Gu4RzqWuqo4iG4UC3dnEqj/HN+odmpGthcIiWH
AUe2V7GlDbl8ASDwxQhUL0kpExVkD3jklPcOyozB7JqrNHSJmxmDuXtCmXhm4hGokRdj74OcUWQs
TPuONPFzPUF+Wf6uuHv7ujUyKGhFNAgnU9WHac8YTKjMHKpMhsdl6PjMg+glKvm5hyt6wfyS5lrI
7omh6iwIQM6GOIMjXGqIajPECUcnteTXV31Tm0qZogyp5tmU7ZyyW2ZBuhR1a1oyjytjUIfMmcVB
Okagerf5gZwL3OKxL3GxUc64bBETRlw4ccGNFtr3UeMFMypI+296QtS8r0MVZqRJAjMfn5oEHK8a
OpaHLN76QH30jQ7tezj9B0Cl+2AZngwtYcOBPReDE1RxpUd/k7osHOPVXbBo6LkUE91W3pElQ7i0
JCQNOr0wYQoKbmOgN7SsuTExpDeqwuGF9bq6UKAAgcbnHr+Rp1mo2s4xzHB7oJBR+6HjH4D/Ix7/
Ae5d1X2ouPJfRNWhP+N9xBY/MjHQk3DMQCLH7RcJRBNQwj7TvDO/dzOe8z9mHZWjCD2BGckMfqn6
OlNc/alOfnPkbmzZU3zxO2aP9NjrCb8c8v00UKt9fg4sGk7soorUo8Al027983PfziL1CcUPF6Tf
yMRomMpfcxQ74kG9fonm5VY2nrs8qe1oyxB0bTIqFHZrzgpTBd8azoh0liBKQSCb2GyFe9SWqlEQ
DSOPK0/DTCLTflZ/+vfzOTwS32br18wnkmWBVYIM+MBzRHpiI85LktwvAGYaig80n8xhB0ixiisR
tGJMXsU/TsEYkFzz7WqJmeUmRsfiueE8QOVX5UqvjTu6qbTX6RJe0PddboX5yW4+ldpelmagWvHr
HmsN7yP7flEyd4/+J7n50bZgXQJnGlq+TJsvM7AH4HfXoSWC8K5hC/AOYTeHaoKauHl85WZIb0QB
vp9vIlW40dKyPnIDqlF/2xkz0gmVzYhl7wSFeVTBoiwUhsnl4Gt3cCZ/WYjH9eFQV/O+gFUOTldE
fbvGPpiHpgJ3fCECr10T8QvNfXh5IeE3dX6SmxrO8odXQ1eFoQNtX9g4KWA99Ass3uztiBh9H/pm
Yr8TPLdm2//iggCUxOOYbmdsL0M6CrCJTmHQBQdBjA3fX0pxQVjohv1RAiTiqFfuRrrnVJzX5AXg
VJMF3HF1jTLdRU8wrRnhhaJCu5CgbcotCHk3fT5s4Cwhsa3yLm/EZzcEorM7cn0Y9blGLPp5ZPPV
Z2QIcb4ASKQn9e4a5PgnyCKtHvJ7eDwZWXbd6BuzEuXVzvRNdRPnYYk5Z2RkbaSzEyra/zpbrsnk
dde6HjQQ8QrEJSUQ2xi7FSW/4mv2KvzmnXsIKvui3rgbk12kRkOCzIf2nOE1hAcrJMfbiW9vShEg
kLGU+z9C8Eo8rKhun2HQmnrQZMAexvKAWZHy1mEfNpdZsrDP4UnluElcZjtzC/MwjC2YfDMvRV8b
abqDEtcZ/l2K/oE1yKauCz/hP6lyvVRZQ3v78+/ixtfi4xRmkIcmagJ6zTpdIqI0FYFwE3jcSOsn
CqOpl9ui+kzeVVZcsPQHgPcCofTBn7KoWiaThJupH+TlvSynQKSoX1P516EY3pYbKB4oTYRW4CYY
I6MMa+Rh+b+5I4hxvCSI3i+iwmkUsCFnBK0eY94z9YMxpiopRo540Ur8scrVtnjg31aHTak8MSIv
VF8kvLxlEWd22lUnVfLrAxJUSipf9xyK4yD7bs+WRlcsF8jNfejkiQfzANnQIbosNLkjxF/3ovFH
/hDof/GckVWYsXSHAzesbF/SkWtfmFaxayI/ipy7m9188mPckc5JqqZohyrCo9mK6cJGyqfKwKxQ
WjHg79KAsQ2p+3KGr/zhN5vzFQR7+yIhR8iy9xvN6rcKeKp0MFC7px2L9TViK0fq2wF3yJlYGRG5
To8wc9Ol2xGcQD42hygxqA3omzS8Wn9EY5d7dksLG3WlhIx0a0RFF3rFBCEoUKAqWmhbQ7ho9MMw
VvZ4eJej95HiLi9wRlrfNEHxYUz5qsor4dVT6DrH8FtnA3Yh/FmxKaJU1YEjkaioE0gACi/hsi8x
C+Fq4H9AYxEtsV92rLureFimQpM0pQJmkdatSczp8LqYQrDqbixnaC/OhJX2y7H7VbvTkUbcRBlw
GEUpqSDZfelS2U9ShSfwuyUsIU5lRwhz/RSN4hdUmZ7NepQyGFt9KUXnZGQO+Mu1QxJlAFjrb5nK
W5qsbpoT3v9bYJubbQVagogoPQXl4yJOEUxH2rqkhwTkkFTenftdluXl2ZebquItF39jxzXFWNtM
kbmNtYsEwHn3012nOvA2cB/VK8LUAMKlKdOaqWSG165GiCyU2PZZHNc6oGuMFaOO6zz7+SSca0tA
4aYkZahy93nmdBWGSIScpMj7ts5hWUoetG9+ch6MBrIiJnBMnZ2SWop9gatvb/9EMZkqoEixmOlE
aq8aqzqDTvo7p3eFEPt+wnDiucidoRap6An5w3vmKfhL64WpQAeTSBNUl37Ako3dYEJtkP58hR4i
qrCr2NIZl632X5MIZQJmmk/6jLoZSBn32Ml5dRBxseeCOfOOfZCGOq4/LrahncjSuSmiT76fua3N
4azGfJQ/43k+fuGtQnHibt5HYEhY1F35xPsYCkVJnIZNFnzdtCf2Ms/aPuiIwX/Yz+JJs0ttZX8K
TNHUuHs5ukwVCfNktKcYEEohwIlBdLuLSKWyIg6xndyeqI4flDXg+92aBkyZO9rK8aM+S2PSsFoX
6B32NjgV8pZ+8qyFbUS8ql/XjVhiyFXGiaGHT9H9WfG0csv2V0GNBjaC3DyLplpBN5huAleXGIcA
dGyQRfA9rWgfxQ5vjzR2Gg4Hixv1svSpx4Mxeon2b1w7bHpfzqmjFao4OcEbGRNt5GvsoXwi0IGf
lwjDTd/yauZhD0M3e0eAOVclNbEABltU7Jzxw+sNwULVkg4MHoqwed/DfbchV3665LDP4rgb/wEK
ujGUrr7bMpK62UpFLW4mfSE/JsA2JLKXGONveJYwlHfV2aQHG43ug//A29Vc4xamHc6/q4M36ZE9
8IF7H5mdLg0XthJImyrwpeXo+WQ2EmkfjOAJOhbaz64SRHTE1v8B/kb2O9W0BShniDxPyPNYZ+fu
xzmTgG2/DDaFEjdxS6z2QeiIT0tfhmxzTH6gerxOqQprjP90GNPz60xqhBNt9DqCkraskpVIH3Dr
FOXYRXJr1Zla4/OpvvhSqEe8JCw9l31Eq614ZKHSV8UfFlO+j929xA1+MCrqEF5azT8iLn4S12qu
pKDBsehNRrz7bP+7ofuE3+rmpEDS5odAOrR1p/mzHmVQmBbjbVxeVcTJk7rVjIBBvxpFpZrtfS9J
CWXE5dJRRXwhVvWtCAcNvWASfc0jZsvFpXH0hQqEaVbxpx7JKPr1voC/DTRiGMAAjmtDJJAjrEU/
6H+cY9Ceb+XEsL4r+Yuqn4n08mwDdggctALWGeWSY08oLxMRQS0O7opWLZgcFDTxa5byo8yf1lTt
+SrPWZksWxbvbKgxUjwF01ayFHrBIaynYasN1vplnB2YBvXq37CcosIrHsvFv3+TK0Qephltf4K9
Y5pjR1ZT9n3pVMPXn2jZOqYOyvmcSZV37DkUszNQSDERpLOKzk2d7hj18IboH1P4nL+UFFzh69R/
SFlr9MRkr8EI74N5H17NbT1yKFv3OmUoKo7GpQ0OhRkMx/hifQUK91aX/G0aOar07mGqMGOx10Uf
FpVXRlgwmyKpT1E+armoNKy8mIUKaxRlBtkmgydzH9FmYudFUM11QSE8c0lrruMibigFb0Iv+8uF
cqrawGJDw/9l+6WmBHhH26YyPJH/8VBhE8WX8I5VPkhPn/8m1fGRt6C6UON70/FBjw0TgfSHHwPC
6Dn7vcWDvVbbOUjZF2cXopmflIdQaR5YGRqzBcebRJieniuHdeUZOSFhy68NAQm5SVLm/gYIoVUZ
tjR1Sn8dZ57pZd5I5Cw/gVnO+qooqZBOmBd0vgB9qSjZiIBBHjOQNfpY+DyIVUH4T7c2iWmaVQIL
95bu1ZAfwHolNXnpyxmQlqZC2tA0sRSHSkNmDi7xry4CzZsTXwUiMsFuoR8Tj5yTPKKoSqcwqlFV
v4LsJ1tqCzbn5P5aexh6mONyQUppNhhtG45JvcQjGKoAA2vzAbiKgmQkL+fNRe7QsrfJRFVUpk9K
V3V2+ARVfNGIHCUJSqIxrnqkHar1EJHDEXWh/gzYy27lj3o25ZTAiomBEOx+ZD/0WxtO4NIweA0C
WMQFxsRb0lPx8ylkoqrbn8Ik8oenxemBZmdIL+ryeuRgmGDFW9s6WKhLzSZHcjA9b99zXVAIjo/e
CcxNqPnuWKfD+flKuISwWFgxVdIcVW2Z+fEaPBpooe8kcdq97oAlo9QsrKpqx9FhfzuC/BX9kM8a
grsTLSs+M23s2RlCqg1GwJK8ifZpVVewV1TiYQ1KO1P0Iw39frmbUHYOMiJGtk+HHw4NVF3i+OmT
VZFmvyjg2tc8zSYbM79741bvbwLjyXYpVoJ1BNswZL1RRXvmLYOl7K9yjtqq/gBNTHtlwQ9A2T5q
Cw+Q+WuXWcGpa2xv3fClGojdHxzUy2v2WVckqWXb1+GS4GOz0ORbrrgKksNawGBhPyeTCasepHa2
vw4yj5UWccnZKoHiKChWEJBcf1EwPwEWd00zLtOrkXzyDB9VHf8z/mhegt6Pi7G1GovHyIUiyj30
kuZoePi+SW5UkDOsztvgGmJUrwRA0VfjCjQxa6/W/bhxAnxkKf2/ceWS7A9abVCSD3HKv8YG5FaL
G2K9q9qy2oRLyBquBfRDuFFd4cO9Uc5V9RYHDVRD0mwVNWWyyvwqPzjpD9bP44iq5RIKqiCxLsPo
yMG5wFUP1C9NSL6wA8qvw3XjGnZGWjlu2I9XM8TkrdSGXZAi9VeaYXY+GeGhXZxrHDGl4k2YyWK1
PyFjyST6ODsdG0VykqV8GkFUALdXZksRonpC+n6ImA1x9MKzTFSt5hmIpvzeoLALSsc3lTyR0p1e
8OCQvAgmDs2wU1LGnlM1/qn5C3jHJA2Lj1/BssCuxiEguqdcDbGH3Jh0z2vyT1Js07L3UP6gteaK
4nN1ZsoPxX2wUU/4DsnEdz666k6eGHEVBjzHDkyinHemZxCfuQKLU46SYp5C8PkK
`pragma protect end_protected
