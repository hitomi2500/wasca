// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aMYGBhRHOYo3hhwWDdWsgGbJR6CnFS1atTVwmKbksarTAR4Wl2fvEd7AhxCwxrpdCbxGTEZkZ1sp
yQ7bgkV0adnuZ002y+l7UCd0sE05BsYvGJuMGYfY2+t7pIjcaRoLAeEzsOhmbyMZ0YaC/KXjax82
3gFhb68Ela43cr3C/DgjhAq3LillLKwzDUDY1aD+ozQ4rq6XZqHhbukUGNi7wVPIKrftPEJkrHnI
LjnR4UtmO7VFONkrhm4y/1M7wZeeIiDlR4fMx4RYH77Y3DXjb8XDxpfdAbcZEZ0MNLzi6Mfvz2ko
anjZ8fy5nlbpLdYVr108lPactIgGAasirHvdBA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rAappjwhmKuW2P+aPiyWs7763yB7jp6iqdmaPYorRklKSij3dhxqepsdgD9HO/DAfNlMbcGf2mNR
4NF8Sd6Y1uav1pWyIQa8NHBSuyhdQHTEAmdax98KusvEUVFjP8+LgSU40u4XXWAS6X7pjszM9XJy
azpf7XUfePk3swTK2tgZs4MFvhFJOge5X6ap9pwg1v+XvModWKiPw7UYss9RHBxiNGZ86Od1Fij7
w6Caxu5KYCxtLfd9x6vZ9EPbFfa/UqEGdPNKkAQtwn54dJSWzsXnMLK7+1chIbfx3A52NkVQwHyd
JOozqup7V1OjHLsTdgfCuZ+bNd7iNUpIvZp75uayntv5iq85SrgJC+JgFRleEWeU8PZ6VYtgG79D
Bs7tFzdCgzxylgSdFihUIGynE2BBWBsJe0IXX574+E0WbD59iaORgItsZTpkI0NDI1nc+ZFuRRLz
S04mY40rV4j9ptfqxMtTbp/i31OKafqOfN+85TdCXfSN7wEnr27bpTerdr55eVAIjbxQewTyMSgB
VtTIyN2+5pfQ8uJtN2y9aTGw3iobDVCaIn6QV5DaYgoJQzOFZPvaezPLstKr+apdjPX9sK0O0j6a
eADaXHRggct3qk4lqxoOk6heY6FU2VK0Cy3bFiVaQAFPLzkEsb9iU7YionMnZwUa0V5WPKiOXZx2
qKvP+vTOPQsByGvSSgLsJxs22+mN61xW00WmEKoI/YGYSVhvfNXnetIKRpeX3XQzjoGS0W3znDks
q8W9eEhhIvYnzP0hbfoTZ01QsJR9WgT5uuhMcP5fXiMwZCDFw+/3y2bexNmVR1/Vt2FXwv+GOIGT
lIu3j1QwPdNUVx038qBQQAvZMNRhR/jMVeHWiTkS++3OypuCQcueRPMxBlfRjQtVRjfz8no/DCAg
yR2irTaXqCkwNtmYnTx6xAKUMXCAK7/fOiboYfK+kuuaf8kEdWGr4XDkzf0gR+aRDCOyx52KN20V
HG9YlIcbki51dLB91LgxIMNhkMkKOkvWOxuE2t3hUSFTgsEcgW/p5SZbJPO6ZomMCQzoDKS6cZtT
PbWiGr7vJ1xWKJht/7zhIe7xzBV6/G/3kDnzC00yVaq3BuaFa0HhReUpiOUT7AksHiRiA8w2KKNX
t98G2Bst7XK1wjEhKfL2gR7aW/h4Q5o4ApYEMwOEHWIur+N2B5zlO1RJdNoIpwp+8/syQ7NS2c91
0lHWLzhO49Ak+JWss1VXzEtZV0lRunMbIFMEcEsE4XN2yK7k0s0WOoYwYh4dSQOEl+Kvfkf68Jl9
cRrfasKYpW6uROKHdSn6PpC2p4ZhprXBgutKI37InwxECeaby3iM431XtEVF/BfSeV/sa9KbtXJ6
V3XkJs4sdJqrVnvcDBntdFqCsyMfkxtfDF4JF0Ch7EGz2oIiOJgvhtAWqiPsbXAdstyLy6c4ofKM
S/IwVyFEz3t8H0bSdEN3+5yEyIHR97nb0+4c/VviftZhrQoCxVscfe+zimBQNcLi9Vq3vSXSMsMM
FV/OwNt8lJakWCXeE/cnvmOj90AIwClN2+YpbI19RrnQ8/2ii8dkol84stJbBNxeWClq+V5JhwWB
T3oeQpeBDjQkWmGTLQmEFbUoM9k2JJoEbjOecnUoHTZBx4MUG+otTtvU0SUMBXBjQFhjDXcsXcLa
ZSp84oyC/ZqSkgaxMTIFe52ofJns6s5JH+fFXXFs2iwbITYfhhFGttWvubqqgrzAUDmHchejp5ZA
pm+3qA6d3Bc8TeN0fnMsg71D/dbGfS0HKprkVawK5l3dz0VlaJCwMFhwpX5V0qARUkCANQAI7Uvm
nBuwd0ZeGFhhngVKw8Eu7w1spvU0e6nDNa1CT9GaJ8S0CyH4z9yBrdT/fA3JJCD0821tMuLPBRr4
nXM+mpPdOLj3ZcUUFzxYHZ3BgZ/HXDdCWfyidqhE9/cuC7LtOcbHcBWu1ilA1mjEU90zDQEyVKRb
u4DKhK9zzrAQG8zconHgjbAnz4Y2hgc34M5HlIZ88b+ZShOizHkXqkGytA+2HIxFRuqdoexn1WMv
xzVGIzNipMzy1ZUvaRbLXxSHkaidw2J2pgNwLK1Sz7DNkGFxox2VebdHzco36xfWHFFB5Ae1VKig
V/EV44T3GU9ZROFVyAA2iyN2fMTIuTzweTMc8ypsEIBavmI51W37Q3ngwjEIK4Z4twmQ5hclQ4gL
6JFVf+sDVFf8KzwL9n0k8SBMYF7qVM+sEgG79VvUiYUwj5xwJ8Y+UqM07iAmkaibNDVAQdAdh5Lt
tCEidEwnMGFSyyW43+JyjyF9DEObqNXxulPWVvCEyfhr336AJWRot+ORHjdayZ2PUIT2JTEbfmbN
7+hNqbcilG5ZA/Hd7ugMQhXCrFSzNJ7kuvTQEpNrffVazwHWNuU4IaogtAV9G1zmZBvMnrQdx2QT
nrmvokj6gXJw4VcmdTV2hYnA9lxRGgKTVFSOE+Gefn9RA5VRRQuVzFd/0C66SG46Dnfnxjog8Wcu
RiZWJqSjKP0swGYZWKMRwAAxuxjenr+L9queFGsjzeZmCFlIr0JFNyo7Aqv79/09ltRAPbv9TxEz
0CFoFEaYcSMw2HVa38Td81YFgcMdL+F5YEeNfT5IZW+T4E9OBfk+rMf7owkeS+QNC4Dktiig8eYh
5GZeGT5V0WKwqf6tvx9aEas7pQJRNUvgveooygp53MSGMKKfOW11M+Bwtuw5Vh6TSXiBSatWLDXK
KX2MBHaPOVtSJsOmzB/tYbemFBccgGznNGrO3dZC+pZtwe11P+QW94iiTAoAvvjAD3B5pUeUMCnw
Z/EwJ59vrVgEUovVDweJdJXHSKm7f5xoBithwRnYX0MT9eMO0ILIMywyX/hpYvvm9/bXPiZfqV5l
2HXQevUpuOc2hRgBhmzc7ZpMBcY71z7oief4R/SeLMAN9hlB89jm+NbTcYP7oGmrCsOPMhpaXDkS
kNlIQ6IKoHAPdMZPOU8KV+GDY0iH8syDN/yGh8q00dJqaGZHAXy8fMWOl0XVvVk8KoV9druNPgsR
PAbXxx2PoZXgEwd26pU0CBmwHTWw+EuzSQMu4uHSmxX9snF/72ZwbVQPBA2O6iFyDJLZapgqkkbq
KtRZNbEB/VQkH7NmetEQg/NG8bbfVFzkOPdq4lfZBnJ8+l9q/HFWxID7+IsVZGN5qaQeHgqn3qyF
2uuQ21alyIu7z6I92w2n6rUbk4FsbKCL8C+K9/3TF4rYA7KwSbvLKzFa+2gYmbHMukY1+EXbCS1s
1uP7XpT4dD8vS/0Taf+/BPO9pjJHDzBeKeUD+pRiN67WiIK8rKREbauBG0FrJsh6saAqIOdzEmKD
6n1jtcDix8uRjzGgkHQYqaqW+y8/lVYD+ansIQchUbxHTFHPXyHGcTfLmA2XrsKNgh7TvyrgZ12Z
QdzJxWow2qL7vWI2uKS1yh6KzzD4MbPJQTeDtQQ2pbJUZv4BOZrKIk787n4CXi2Z8WulPU1QdvUi
8ONsSjgxeKKkAnrsDqxOvxhWhkNOQk/DhvNC2UN5CkWvA8MxKKLMI4bev+76ET39m1ZIlE7nCfwt
eCKjRvc4a37CFcpaxpuVYSNkHM+52VJKvivP43cFsQQlAIJEPq6ApmUTQfKVL3rPMqdes/WmQji0
OjKFpxEp25Zfn1IEWRNyRk75WbkoiRslnmVD2ycyQUxMeUj/rseNanrYUAjbsz5bJcwusG7t8cOP
kJCTEmsRcmUP11hL+m+gz+VnLCQyVljmU52Cpu3pP6fslvL4Nj0V7fME7cAOavhYf6TW1U1ST7Bv
4VmHGSVN9IsvFVTnfjL1ZIVuAo7IAlIv12Y89+N4FL+CVBjuSbMZCKELGh5vbLSSmJjsWQIJvXuZ
fi+q8I5KyiQaxnJpMQyU1JJg2ERn5cuj+AKN25/CPl3Ad5R2GXly5I9ubTY6Abw4shWwjf5WQEsZ
uTA/876hNFsl6f1WOc/xq0mqx+rm0Gs9ZPfuIYAjvl5t1zDDT+sCq5h8PKOr9XYHRiRc5rSuhUmb
WZv1s48yqbZRu7olo4yoDB9SPjHuqp5fsNhiypWhLoKlnpqGnTlAPQ9+WyMJUmbm3vic53LfdqxL
JPmVTkHL7BAiIx+DNaXaypC8wQf6eeR/QuGDGmYcoWPFwF5WeSLtxhEQ7sKGWfnU4csIA7AXC/dR
4+u38/8TmSJUZMkm5yDeBA+JkwXg+t3fOR44/MQM/7rMQFY63YVOCuVBAmPL6YF0tKwdLJjsJ5N6
n5sJ27/CPfaTKPV6NZyfnKIjC1bmHedi+9aXv29XNFU+4KUWK8DRTfLhpmWL6EIjV0eBLSDZ9gaQ
CVJMWljuXYvrJURvDI49F0/LdL9DK7FMaVezgY5N3VACekYkNXpb8YCpbaiN+SncVR64d2WSABfQ
r2Ag3E+nblt3NSqhSQC1ubwQuf+ogXB3YUHYKVKh29gNh2KMnCvsi5PRPCWrXn7aLrqy2zgvMI7S
ZiyuauNUa5fJDOBI/y6y8VM6y7HYg1ILwD4jv12OcYRIEqIRdjJotm7z2qne3HMuQXovNCnNkvo8
tFThcaeAdWMBKCSS03WzoHiSBQvDu1tKtD5hXCxfkUEN3pIm8LfJUirv6Sw5vZALA0jpwcz1fPMG
McVe/XDBwBdslFX9/yTLCb85nloUDxfzF3uhZcyh+VbNMTL2aYKHPAoJEF7Kw3omcUGUIWxk+fjq
lZSYjNlRKYosD9lNMM8Jhh+Aa2gKs8/kMAVY8uEpS6b9obys47wFnPsy0szkIavT/TJmbRDpD0ta
gFIel61i2w7xDNnq+NWx8F01ihqYh8Q7C7RqJRS9k/zsnYPORG5kjaLTEa1N/NAilaWv2y9h3EQK
cnjzHRO1ejXErnOxqVd9kR6Yu2xAOBUbDvUwGg75b4Noo6KMEPZt+Ux2mtceznZ0NF0yTGqwn4w/
NfG3IhjQlm6sOHXX1Z6gzuiFBDJjuz2sbm+s1pM0Gn10LwPp5At+aXlConquA3ZzG/WCEtQEYsJx
3yFdMtngHJ8IFmYN58zJT2nDPOcCtmoMaDj9y+Ykk8G3sGMnCqBlo/J555LRfeQU2wpBTE76I/8J
uJWLY7y6XMQzn1V6l5wFNAsEsOVwL8LbIMR4h5W2bkrSzjZgUZGwFTkTzjsFuhTVqW8XZXHJT3LK
cNamSRo0PnotHRy9MeOSp/zW1aXe5qrdANqDhlflWkJrHlBCV/saHBKLOBSgeE1K3GCeX+ZlkVqC
QC31+kVqEfsnxu8in8rP34fQT4Dbq5MMCsIibGqxVkmPVDYQFLEj4SB2vNa2b/L+4SZHQ7bkl8rE
GbIpZsIQt1mOOJHqK3ZpB40g6mdFZVYGPhRtJCc5xkb+Fl6fbXLA8OjLpXZ3v7MkRewn4qXQShDS
gjZsyTFalGwDKoRUUDTHRsU2LpVR1UycyP9dnpkxmVGeHaFowAiHYxAVv4Cg78V5DFncK7pG+8Cd
pTEne+UWJWvDDImzcLWaBk3nSUn1R84Wv+1M3ghQtZ+ZoWUqAOJkBKyB/83OxTHEH+QTVMzhAgby
HCqtmHK4VC8mjwA2zhlvvT5Yyy0gg2DYzngECfMwh57IQEsitqtXy5pAhGIi5KagSgTjarzrLwqM
nzJeFaGYNkxLCPHeeaaG826mR7oTcwlA5rSy45HsVXnJ2RwNvtlaipqJizYbRqH8+mJFZ4LKNPZp
Xk/rZnXua0aWzI7643RZEADWe38TGokikcH9CgEvL68WktxJnhSSEcWeyba5f3HeC7rInPA6aGnx
vFZQIy/PAcmNq8gagsK0KwXw3rJWdEimho7OA05oVoZ5odGP7O1cauMNic+bAHy8UnYOPRUV8IlR
+eMHJUbpUDU6gbVMjcjZs72rNxjS+OwDcPp5OiRcr+Nls+//5HOYawJqVQCK6DpK8b7L7+8Y0A2j
vY4uth8JdsW9IfPXoM0LJOEoavTckKPA8KZgXdyre4OjrxdJ4Hj+YT7nCo/vc3zoOLezUmqTpJhr
KARKAbauOfg0T7CCwX+tWJ6x7E28g3dmsyUO9TXpPmdCmW6CagBal12bpUCmRjNVy4+phi+0b5df
iSLk0dBzn7c7nulchKBuo01YT7UJFubHLFoxvK6tLvRK4l0NI9yww/ujoy2+6Vzy2nEXlKK05Qyn
9grrpwRby7UfPJfeA1/ARgfIj1DrX2Br60k/TiNAU7O3gJ1JOZ2csk6UOwbIypoInLAPIaQiBmAI
aQVgsrcbspRaYugWeFcagTaRNyatHlS9q0A/ci7GKrPSIVqQkPekr34rU+7pIyr+Cy3G3JfFs9Rw
dMMsUaB49UUAAv9dXlZx52wf/y8domUrceRcZegAuZMk9RDldJSpnSpwhqYmM2+8alEdSNllLHGg
MU4abyTLXQ+zBR56/nXlSZo/OtSDv3nyiMfJUjXPdI6uNKydZxntFZzaRIA/ULfY4cVCyr+MGlEj
1tUS0NXmjP7e/in80lYPaVJeYFfjmss/CT9t/+M3bLsiAPlhl49X+hSmyYXYoYMT2RnrKB8cp75y
lskwKBA3V875JI6yj0QzBIhMg4zpWrb/d83P9HH36+iQqen+1EFtu0x3uY1UnAzjpeBF/8FZHgEk
ehvo8sE0iS1YDK+ygnjbRG1KV8uDL85DEMxQXd/0hGBi+yDXd9JTW+At0XJ2f13KmGdD2U16lnMU
E6163/WBfYYpZpInXZQzVoEtv/mFrPfQU+IjJcaQpVEbotbY0Dh04sAeuI83d61svlZl6oBFbSQR
g/SLxQouy8NRGeG6fyfxT9n95eBOFwZOT9y1t83O/e3NW3Mcfr517max188KEaH9gvJmrwRmHiBW
CB07tt2xGuxFdD26njlzyfWT4MLH0zYGhG30KCFJ1ebx5MB7IOtMTZsmCZxKNEzyikYVJFWW90sL
ia7t2VrrW78mxmrQ4MNb6GeLpA4ZADvWU+7nmIlco8tvL4d67IMtYOdgmvKvRAAAvg7ot767QG44
4Xzf+OuAALZM+uDb8QinUvF0Zd9xHNajldmdffrTvvwXHVPD68Ftc+Nj3+787HcjSAuGMMb+6HSR
8YCW178wc/SM1F1S4VCTI9Hw1QDskq7XSAYZYuuV6x6nwlhR4Egym02aW3VpX+R/3WoQ70KSvPC2
G0RRfudlGe7JXAUFfRxooUNv/jRGaRaHQcOydSo9iR/w8Lv16LRHWD/eNLcOXciy9Cmf23IsEapU
IMaMjihQKD6w/X1yQif5+X5oJ88NaZOk0o2XdDsXuPJT/i9KH/Usv4fWCxzjGCISk1XMHrLIW9oT
6mDrM7MauN9ED3iIKQgF+A==
`pragma protect end_protected
