// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:43:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ix9FXWvdOdH6td9NnhiYLFWquBtYMQGf4a+qPWj63KayrMbzXGr6s2Ng7IfYa63B
ABoFJNdTK2piy8leYMu7hbp3bON/DTIx+c7GF5vJkclD/OlBwPn1GVfWeryodvXC
FN3jwx9QmlYaxsUXQj6OFTO4zBz1/J1F6xENsVCiULY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20672)
xv+5bndE2YC432s953C+jRo35NovxjzRn2JUgyCgzNbt8XXTmwYvtVtCGz5jh6EC
EHF0JJRhAhgDT4Ol76xTCfzjs9vFzLxpEelrec7QTvYFVmsYzbZ8Afy1G8WffLFP
7N+QQoJyI1Mx7buuIbmh4WCHvX1aC5AeJFtzxOVKsfc93wRVw4Kvw9qNWjdVcodH
KtgJMF1CtmRgk5BjZgscGJwhkZYAwuFcqv7Qwo++0GaKbR4O/dro/8MkEewoo+S4
0EYEr7PlnZD+jCbIlZLCVT1/gAP30oPeswZbCwQVYsDK1Vnjpm34FdbFjjUDiB9R
2FS0U2TgfEszlo7mrTVRSk1P6nYunqfVgMVBQhNWR8JMNDuF3zWnSDm8owejsQH9
5lsPORaYYPerPPK8kPDSH9Sv3bxK7e/iIGoosT4gasDxdjS/MpP/FQ8hzniO1gkr
+6MLrt3VNAV8If3aYfKQO9M3XsIoAKt3fVe8bifaQeYQ9FrkYU298sFXgFabnnJD
Two5qIrTsO/sBeHhaiSRWs25dvgx6cEeRtGduvrUe1HTTHSeMCBXTdACVG2XOTN9
h+85b/nIrqvuTWTZaY3mzuXxBM7YDbGHstH0LfVFKVh5tQsz5dfseJBIjWVKBQdL
9O/gwsziBSYaK6hoYrKc7Kxo6VlFyHzislf37WQdDK7Wkkc6vZjdM/6ABwp1eXzw
+ed0LvLDlkHKB/FmnQohD9uP+BePhZ+IfbfDrBeE7xrruK4TvDQkhMBnLWtqedtn
a0Hqma8+wj4EPaOc3gG3mIrGb8G96MD6fmt+lvJdZHL0Qw0s7E0pcCuQf+igR3t0
hxluzvF5qyE8LfGZFLraxoEf6R9JPcNYfUgtCz+H5Z7uGD3OZ6sQ2MidJ2QGsCO+
zAFwvXDN+EOOgdEZZdlSXRxKn/Y6B8BGUievlsN17cvzM2hdLDQnNu8vYAWsDyNu
uftxpd20NNTKoT5CPpMT8dk3jpvDeuYPmd+GsC99csBN/PG+GrhWRMsbEixQW9bt
85NxHfm1ob5n93vWwJXVVvzYlD6XxRRytKOUFfx+SRmEzl1+vgyuQnIHOdRE8V3x
SMiaaW1nGtPpTaRLDoRo/rpkj07Vq0+K0rqDYz+He7Qtr8/3fmMV6Ss31WzmKpag
PqEMr2jXBHqo3K6wyoZwl/2fj1SoB90pS8cY0/SBRW4mz6a4MhR2Va0ErFRowsI1
dFwoDCEuJbrEhF+U/wsOiNNbrnNF0f0cKIsy0Xh7GesgIxd0sCn+57SFZ/IvE92t
G54FZ8XeeJ3LZEBmZUBqNJCAw6BgGcCv8CvVtzexlY/m+3hdZPvicgOLgW71GqBU
iI2SHmtPIgcJNSCbQp45yswyhcVK/lYoK3oA3x2QZYppTCysKJMq14Uu3fTMu3Mu
p5RSorD7ACbvKz0tviS+OG63qV7qvqz0Mp8mmmPB0mR/HM9/2bUgKu1u16vTBhU6
CgACuzXRZxEj6XTaozAfhqB/s4BkP+E/USfrd09zryKyxt6p25MT1qhJhMvhIGMW
8m4CsoGe1NQkHZdjZ6I1sIp+KsJ10JXvFXg5bYL7XP5t6U5utQOlk1wzfM/Xuika
LJO/Xa22XYFDIPzVk+qUmFjeY1L/lpVh7AVEv/zrygSSkxpqwp4A2bQvMNh+lQai
n5jJrZueL+fU+Twk46AudIzH4WymwcwpYxgqZ/snnP/v7Qrh2Z1mVJKDsJqeB8P3
Ol+2kSs+PtZ++f+qMYycVqXXgSRz9xfQFh01GYcGn8d/mMGSGBxYEvCbXdE9Xtmm
gneg4C+jMFQChm/o1V++lE5jZPgKUsYBWDnF57z5g43BCSlxqak4ilTL/2d8B2HX
vAMm/GVrMJOAElgWPEbmXH5FRJrQNLntawNqgFJ45YCKa0Q2qQB5fRA378bBYDei
rdOuewMTBT0e7fJL4NPmHlGG8qpWu1WAd0fWJ8c42KgYyK38+Us1sU30Kf6rMJpe
3XF3Ld1lNb62cAhP12LHod+G1GREooUuqfvLxI8Z5piDOv6s0xjWjH3wzoaBpKSt
htFe87m/qLNtLgMsh8S+MIaQllDbnCzNQmB7GnlJBPLUoNvGYJRoyr438Z6RefAW
Jq7MuWRZFDDGvryUv6xQsb5jQxNAOIf25jAe5YB1XjybHHWjGjJ8m6Y+Cx0ZU5wr
EC61Fwsd+47rt+ZsSjYVAYH4AKiFdSR5S5qw74rcVOIed/uN+waOaN/XbO6DeZvn
ixt45UJEXWJdM6+pax8OObqPEEHEaUsP/yvGwho3397aTu3i33Z9hEnW2Q+04m0/
Rk2OmJIcLla6fCK3jBdLFGg6S5h5MB6MAVvYiu2pawfE/3JYmmDAQUz4f573uHjC
2vkMKTHWi/EZJI94cNTbUqc8YKAZ/Vk8RK7JwDtvM2LXIQix1bOwMP/91rpdfVhz
Cp3aJWxBh2xze7kzyKURzPnPIssBLxh5N5IhhxCic4JStIhcJlP/crV1WZqh+Pcu
WOPu5OEX0A9q93YVf3EVZrxGVNCehfqKZkBkDsAGpphQXFPLV0NkV9Kshlm+FKra
aZcwPoAAVZJPDJrf2MGGwWYY1QeC5FLPNcCf0RD9pOHW7UdnJchrv5hslexo62Xz
b5HhRsKMIuKZ8c84L9XN5Z8dLWdAjR7yszndvasiGH0IejJnRmqz7iN/eW+3IPoh
VEraq7e7w+Du9UfxeLe4jvIcFG3ylbSz4hOpJcBX4ldivJNJDXMYkiz488st4h0k
MIYsS/i5BxkrpC0mvhrAamzXveil3oyqNa7QGPphG3ngNFbXKkI69Zu/0pCGFPA0
NSWa9rmqUIXYKVHrMsRDqOkioeDYxykaHZipdHowYYzTZixevBzC89YRdYGrawAX
wpkg/iEsRO91Zk3E4/e1OGNtOvA8/2IRCGE699G7qE819kwYyU6Tzv+EwHnSzQNJ
YIEgtDxw/Zj7TStatbXwm8ui6HtBMwe3kXOIKsl49cjxYGUrxccgtCg+y9C0gKuw
5LbCyU2h/ypeTpo8lJNW4p4pJehC+SG6YYsmVAzabXTQgrGBvVKz52rU6ZKOXljR
hL6NNLXnDiLD9KS2PHhXjMg1c5xQZRCHjsDaRa+JAzMtq1MEjREZxnDj1TBfFulp
sRw5wLgNk7Zhsj5L4Haeg0SwGRvJXDr9yrx5FscSb+9Q5wONv4vYHTp4W6VeKXf9
gdHfvw/C0Uf7+lD4S4B6dJWYtUoiHPsEYOD6Cjo84CcmR/VgQBDTNpO7DekG+YgI
gzLN8ApZrB2qf52GhbeIHWu9RvqnjoXoC2UWB/thXV02waEsDXH1tSqEMss2IdHj
UyrbIhP0wxK/D4fWTdQkQWBDhnL4RCJAd549c0/WOtQcYorNednKW5tRAZNqp547
aq8hA7soomdUp7n5crLYXxZ8lTUmRp7szdeKoVWKPWmaJZl0AlflD0yOfvh/76Wu
vDG/vx9hEvWjsnqZsRnqouSEPyUzV0yxW8JT4x4dtluu2P0a0MewbNLq81oyO0nk
wWfSMHy2/loPID/1P8znIkDdzejtZ/dDH0kvcgXJijOf22dKwlM4+bZUSnY/RoPe
aTapkdszH8BuK9U+zfqcDiTy4+LCweet+KZgeIUbL9Qyae95ucPBOij4Wzv6fdqk
h5yZ8SoGhLtOAHv8saacDfHWmiGg0nKUP2whNfbEeOsYUlhuTxxEVtFJ4SDM/Iwh
GKODlrt9Krl1PfcywfgYrkCP3rnQX7XwTnLqwN1cC9i5Collt/2fCjJLE/6L+3wj
bPKQuJihy1UPABPz3nwL271Niu7Oxhow/0CjMvhzSKNoV5MG5rcMpOwubm0pSHro
vZ8DZXtuispblvcPpLCAeZQ95OaB43ck/EYymiuhPK0dUubbFdb6mVdUlQ2vQPM9
2j/J1NNZIQlZlfhNvBBNDYVvuavRjnQKQXOVYOkDIRo+7/wiee31rLF/XhmqhHUL
bvJTAWPlBxD3Q5r5kpSJVE2IFwkP31J0yBRXHhYh2ntHC5esnR+18xts/P5IJYIw
bo/Zb2lU/X5SMZS22bUOsoZElP79EiNlroocGZFC5IUagOArPdDMvd5aOx2BjRvY
dAQBRJySDs7BGqVD9ad9duyqkSY5/Lv/oO3eRWo6VKtbGU9esl/dsirqb/effJoI
cUkkQC7wUqgX/bz+H6JCGYpfoZz9bQfGmoivga/pwl9e2hnjenf564IS7IoivXRr
sbb1y4y+AZ1k7c+s33wgHjMcM2FTgXZcAdCQf0Q43UPj1i6aJyd0oQn5sUJx3Sg1
LbWpsJOY38dkbHW0T2OuWQ9QRzwrinCfwFb2fW10LVxa/6NRaPl3gY8wUTASq/Nl
q0WcC59MxRWzGRAoCSHYxPRufHVmh9c5EX2PoxQJa8vOhyvqvNvSfW5x8VTNbbt9
cqvh82wGzoRXBoEX2oOD6zHuvMbc6bTGrBSfgl7aH/GFZ8mE9nqeXI2YfhhKIEq9
DmL6Nx7SlNQtLhOHOyZE9wN5XT2Hc65o0Fmldly2IeMd3hxGzSIVHv+bGFYgE96o
2QWMGfU57E8+1SsBW8bGh31OcHAwZ5RkVQ+0nfL1Yr4EJCnCwDGuTbabZUA2HUi6
7VSrvRHyYDnRvDKX/le0sDBwIK3MKIsd4vfTOcNLppDm7F0duiiHH0dMz26Tz0B5
1ozuSCl1hb4esRUqO/jrnpUfNfhRRchJg2cQPTBfX7RA5RjOSWyqRXO8Df3lBvdf
X1ha0rERGThya0nAuFrpmI61c0idvaSbZxNF1HlzeF+JFIwtSY7H90d24unZWLQr
lv6JY6nrRfT0pTMlpPPqNmVYoFWFOcexMK2MK9DZ7Uv7quF2CigpjdzIMzPapUBY
Y+TovAvED8zFhButPKtzRzo6dtYRCNVcRwb+qa5uefTC4DYzPz+nSauUxtGuUFT2
um8eJp/ADIi6VHQr0TOhyJ60wdE8fCmLL2HMYJMQpbGmom1KecKcvupQnz0GxHVK
x0Ovi/gDhxHVUYvHPeHr6LhAJVPWd9LgeAmPDfaTD506Rbip2Bl6RtKRCQ96y/dZ
/T3/LciNwcJvHWGsja2gEN77ly6+mB/95eIwZG3Y8AM+18kbtdt7eFTMulNbBIwa
/rp1dwXIR5W9ohY1epqmjPHMBTDljO9agneaZrNgsdwIq6sWUYjyDgJOfA6b3DJq
9hKsKzGZd9VFbbnm8nV/1Qk2W6hYNbQN74h0rWk6G4MfDe4+ty2d5gT7yo+gC7s9
YLe8U42eJHpkpn7PHJSj9ko3e0kIcp9OHx08fPtr1wvsYf3lbndrLiGOlF17eMSi
9Y+xYRjklpOcOjysyUXeVQmVjAUTTIP1WEVjeBHGFD91BR+85eZf2oKOgqVfEU70
Irco9/BEjSxI5tK7PXq03NSccwwGYlaq8M0gWVTxLCURtVZnC7lRPyy526S6IfPn
Yjkf0k0Q8z3ZGQDyGeRwtUY5Hc4trkl1dZDZO0dGUPRwhNerQoJhkJc/NTwUO1au
KOT0yxht/SqBcaOiI+bnsIeHzoQBOeAo4bbjKSZa06M46fGfNrvuWnEPHs9sytEz
P15ni16K/1a0vmd4RA5DNOlkm6Gqsp8KRWDhEic98AOYFy2tyr7qqVUe/hXwgTaZ
JwSMilbLKQZZpFJKkHHdnHiiITj6ro+wS7c9O8Hsf4D4VS1I+YaLedg4yWsjVkcv
olvOTfsBELcUBF/AScF3Zyg1QpXsYcuGih6hvwKJ3DOiKJf4Xz8yJiCu8Cc1wFlS
xF4ZrhSGBPFYLt24AgXPmZD5L5ap0a/quIjpeilaOaDkWrt6jpzx0Kp4SxyQSVYf
a5ycUXG6jymXxIJKhWKRiVYDFuXA98O/X8jUusEqZ0wt+y1C8zqC+jLriR6HfX39
exyCCwdfU8RcL1AY/6hWpueyB0vltajHKye12iXIMzyrBoct62uj8VbvCufESF7b
BVk26s4yaeXVSiVkpPshblNnMPd+hTzS+55Vf1XFENokulKCjd7hT3YKUr+vBw7s
SSzXP0Zk4SyhVpKbhNzrGAVEcvWC9QR5E3sG0oWU0SGznF/yaIfY02g5jcUFBqV0
UfsPwEf3yWD8RrXW16o+eGWZuokPQu39VSAZ/adp/EtHPVt7sVE7G/FKE/doYi3K
9aHOrG/75nYx+u5m2VOZlG1zdZnFgAa94+bj8fi8G2a5KDUPgJhMYlEz9zso/mvA
ni1Uh+ajj/Zfk8ymiLke3oxAF6Hs7k6Rfh7KV4QGWByQvWsuCPIUVAecrU0N/Pq5
PFpuOcBWRnvbPEF8gC0FvADxae4WJhgTbt2koUmnXvepWDuwmSK3167nQ8rhAaNd
tmGW7cAKFQevQng/RL4/dWE+rfvs6TMWumUXGVNLJJE6zqUEdCrdnQWU7IWXFlM1
hAVNamprHTMy4lVQJ16g02xuGzVfg+7oOv0hR/rXfJAnKfova39yuv23hNRG6h2S
QLPC7prQGbox+5bMrwQtp5CXUTE47PBjr6eMzVbwsoI9/mT13S/i+y0/1JnAmi/7
073wiwxxYYbKZi80Jdc0RAx/tVUvhRWE79Rwx4kEzrEhBNF6sJvPrEzN+oqWrsL6
sqz1nfURemsa8H8rs05ABzVmawX1pGQVj5cq9QLw8A/V9wRn3QJG+5f5uMb76h86
C8A6klFTED0Qg23wrlAIP8q0DeF66GrSJfntAAEo7CvxL/kMlfaRh58qay1jOFuX
K0OUlshwc93ujrZ2LXtjOSeydgAWlFLYtVBrXjs8DWsmCLsDsyj/4ZUDOvjPKyAQ
+LBGVYfjSraN5eNyyA2mFb/GcwEF/lb0+Zd+WKj1x3PddA86mcG0gNcWf25FMsG6
c7bhjVuSbA7LMunVs0PY1LgStDncAMUNXfcqakhTgJDIq+MAA2WN4j/0Y9dYLFxi
/6JmXvh/n8z1pwreid3our17kHTkzuO5+9fwq49aTWmIoHxZu2D4cD4tP8cqj2Q4
MQx/N7XzivHcsnyHQD+N9i21TQ7p7YE0PKBku5XLabL6lf+72CPpUeFRIIjkNlpr
6cXDGdBEwwdIWbxkUi/X9oLu99HqaRmki5OQZwxR2bV9PFpVkC7jkdEjTwqJNbo4
YWTacmV5KGcLdUHUvAoBdgSMKtYM/RdXi/o5JviATxjRUeLW+DPcX55U7OmX19uC
aMXs1tjM/VY1u8UmoGBeDObadiN+31wmi07S0aE801I+TNnLJWWL0Hkk1otW5ru5
IDiZ3bLteISpFk8+LNXhn4S0ynMLRMvRNWDJvnt8Us/yNH5MWjSsH8DIg00o7TRE
FAvebdFNdsWzYNAHlHYUSPCdB7wbefSSdwI34bG4Pr0vz86w2B7omiTzwVEh3njA
SNzt2Ghbc3FzaX84dhtAxP+e1B+7WqIKxZsjQlJuyhM21yr+hSxRy/Ie/7MUsOW2
oJBZ/pOQvQyk2Y0+PrWFU84p3ltzntk2wdCIp8UHo5TV6wdbPLbixDwa+zxCKSbZ
2hjyLRB3tPxEiUChK3L6OMNeXMAXLCNow9S6yByjGCF3poR6ulX9UsWq3BllJrFE
tyf/Mo6Bq0KgEXKCrE9OvTQUZyeIdO0GuIte8dAipBRj8bPTBmzFZKB+sb2xFBEi
bjp4hYnDrKfzcZmv05/F4ED/loQZQudfDTDF1s699NBHyMpgzhVsiQdwE3cF+5wj
TGteccbInyzZ5p+qpWCzrIjwEJQlgfC500qjj+lmbjVUSH6kwZzsTGcjJe/hw412
3/6e2jNOEKjzh6raYaE+jeMl4bKWicx3Ed22hHKZhBQIgN1Q7Ag1jMWnxdGz6moi
3+p4RgYFn7WaxYJLG7kBOLE6jIpAiSZLCcrFFLu/AVD8l3DSSkuEVHt3WBqaJNgm
2goW3BYXIWPW9MB24ZdoOiC2yzq6gyQ3L/FStlwUtNgjlFCcu0kgFNuSWiD26v80
r25fQaPbqkGixoVM6GuBs/QLla6Nd7Ubjii1mwgUK3pVpr2+bd5E2zDX0kUF+i1Z
rDk5Zg7sWP/OqSpO+lcEjzWJTx5OUY8RVRw5J+txvbZXsAH2TZIEq0phedY4VW2P
1brEK1RdXDRqMDlhVTw6FPPa/S+uE2zZdqV/KtzSST9SM2fr4egwlo+nQSHN71be
bGLktvwO/Vz5ikW5UR7Tg4een8l2BGDD/M54O8EDYoKeGbgBK9ZQNrSynG+sk7Ur
6nSMpPDRtgk0YjV6V3jizX2R7CObfGTnDiktHooLefB30jLm5bYxH8QeQlJMbwk6
qa63bVfnXBDwLD9Sj6kXlt49zUPzeBKxMEPXtETZ/T9kOHlXQcn32fnhUcIYYLwm
ygVTR1L32QH5cFLC/9WFLoM47xjQseISXH+K29D4gsPkGdmE7jzgtL/USW/A1x8Z
bUh5u+tv90njQefMuZ4h2LuLbSD14D+T4nUz8LHlIWccj3Zzg+kGgYKICfg9wHOJ
CgtX9OYP9MUwmWMCxAud1cn0sglizsdGeJCY3mOmTJ4LWMGBUy9sIwwDtKBabWJI
Pmvj8L+/AriUBVWFM5kpaSzW91Ojq7/yS3ZTAW1FjEtAt4xV5GwP+a2xaios2sGc
U8OUXxeIPIhJPms4r2f1xJs4KHyraLOvDrVlr86lx8cIphemdolYgEm6NIYRpd2g
Yu7tI184bIPsTOXC1pryoS8MSR4Gqud89EdhmZbFFRQRoZ+Zs1ix0/mp8jrJotpx
f4l/Lh46mcSerskqHXJvTt2fqcYS+GDQiI481mu50uObBRcTx9AkTiDrecoZv1j5
8qNtRvDgdJQLuEMQYvgj8RJbRsKZdxu8snT/S5wxYoILCnMLvjjo5vGHINBjBBeg
+fentRZBkFMhUNX+H2gQ3E5qne4JF8m0WGirc3xAsfJrzuQN5VpxorpCQMHQpts2
6PBhUP16F890jhoAg10dcfdeuP/MsGxtcWbzGLwiEY7PocJNHXyd58vchyyesKrx
8oRUcTj1JnyCGdPYdRGMsgWGx/dPa3r2S9CrrQfatbSQqmZg5jlYswSLtTTlTr6T
9C+THxChhtJI154gs4yGJD9TAdt4sAoKrGISzXocZbGzMdp0NIMvqwmETLo/1lHz
BkHjri5Dheaxpwa9zwjjpdwFXJQ/F6b5NMmARjlsWoa87HOKTbkpPg1Wob7OeE4F
oKO9YRWn0JQET1JXDQZml2Kv1N0XocQ3wfDSVyMHb9TtOdYONzC0IuYqVWzqM73H
nMCNWqnxSTYy71j7qk3M/PBOR2vwxnYbsb2Kims8IGRXwAMicYuk+LUdQ8hAH+Aa
gpgfUQtdx4LOsa7BOZ5FZQYzeZeVA7qFunl+D788CLG6SYEfePanRJsDlZESMU6O
1fhJXAUgV6uWAEhWQth5j5XgauJr0F8jf1OCktQfdHbf0GK3iN2/fCi+dSg+hpQs
d78RMsUFLyVQv1i9K2UMSy3zbb6zDPfPM8d1SS8MRUO+KSW83J1XhagC2oJ6MwHn
ByrJdMt573oiRmG/odGUHT7Rcvh8ZU9egrBpgeNlRrlBQZrNVdCAgbB+bhnKyN9+
DgYveYcyBc9q94z2EvZq5+LZpBc5M5sqryhXAhQWPWMAfoirRXElHXKUDzCc6Xtl
nSJE0dtNNu1pbhYRywYMuVsG/Ycw+DNX6NR8YDmH5gv90bXgB3sn0zw7cEzY228g
dQjHlJLRCmaESOBLkgpe6A5v4uettgovELNrZdJSYKcJyj2vfXOSv7/q7JUH+4fU
8fVpWpDKo2qbqQkTgq6s0ik6o2uru152gd7YSUSXENJxFG7WmeW8Nskr7HoQAl0J
6oGWAKw2GEoPq6F7DHlwA2Bv+5vkRfdN7k6KtpJhD5h+45Su/cdHxSXkxm1vDGOx
ZJIA0Y7TVqz/U9wGMMKNxjXuTuaTHJcOj+dhmqbcEkHWQIanhTPh1EXbheflWo8i
s+5WWLTEKAczvXDTpYHLnZNMmz8W1yDHIF2+KTVVvY4nmTinYNm4u5uDvBaKIT9J
d3aCi317rnYCCmosDSPEi4NtIZ7orSczKIOhk3TdjieFV7HFJKMr9jpOoXkQhI0e
6kwHKVqOZFE+1nZ7cx/+PsuyxlKndPtYS/KU5MPk7cp2K3YFzucz98/qqcshooNo
Ljg310NdSrk2E0YEDs+1JIptCJ3OywfsrL0xrTB2bHVHMjF4ORd4XhgbsS+liMto
/I6lonEw3xBoUWvK2n9tbpNmDcT7EpnJFltfn50NMGNlzbbzNlpN8lsXAGzqz1Fq
hAUXOKWQmr4KsgMJpTLy+pUqaVFYjpUNK6l0ocJkZetFQEGA/LIJ1u6r/SvnxsUi
oyoHbexTRoBQPR6dqonLMa6RCY0bdnLFQKd1NNdBB+XrQWsbrRrue/0s7bR+Uo3E
cnwTdvLuRbj/eGVEc/djaOGmLa8cBSLlEYyNWhi8DAxv27Wbvwv8iXuDs2HQe+eC
+unbXBSgX5KAKU3vo9F8CZftuIgfTzT3nYyohIS8WtCtqTVokxUKtjmFNiU86d/s
6NoHvieY+rqoKIdvyTLPEw3nyGajapLR8UhJ/MgvI4gJpiDqz6NHknV8eIrFAto9
lKGYBE/qRQzmXlh2oHVcwt1KByPWeYWOlFTDxaxymaD/lKZA8CnnUMx9BMU8x9iI
s6GkCnD+1KNLAjQ1kETAHyEI/593nCaoqn506M64EuTyY3ZChEAMCiuqwVnqfTh+
/AoLOYM7NP78g0/EkkfSV5nHm9kIYZu1+XstY/dnEoC/hyW+9lZtmgGV5eD63vfo
sUIFWzShVRPGztOOi9I/ibW4um0dlXkEHv88qP9am9wTUiaS5grhUEurfYy+eKzO
1mnoQBhOAq0VsQWB9DI/W6AMvUoG82G5prNbJ680Cu8CGXuk/AE34wNbxnHW5FIs
Lx3e9f4rdPEaf1zLdM4tf2zIWAMDe9TMnuuiW9WlCfjdbNZSzBiCOkTuIgHtEmbK
AhjTNtP4N6M0AxDc6ZFRI63yY40MNlwDkTTaV/y638neLFcEzGojXDo3pl6bIv8A
yYFxvuYHg0Ne+AtDdAUyI/mI8ozBBqLZne++Ot/qyhpUBO601vCaTULnY0Do5mU9
PuebOPNXWI1mHW+79X3F5tteZLt/D69RYlSnDtQfiu/wStB+rwiTzeo3Zxu63eW3
O1klUtNB+wnsUwMEqyh3OuS7gfbGn1XlxRLlDg9o7BW6BTEPd6SnauBBsw1EIeBf
Dcrb2JzGlJxOThVdnYFfoIVieg6WPwqhxsfJEqaWc//jIUpPJuCt735gAmdsUqcc
ayvOMwKRLqm9nLq9UVPElq8DnM10HaQVyMEULzxTB0Sd7/Idf+6C0+kLgecoeSBm
LBnUghFRLSQ9E3jiS65T45Sj6+HZUeQqQCaAAL8ahrSgha+KrFb9ryTM6zn6FqZT
tgP+hJslZYCO0Ev4dOoFKLzfQi3WYVc90R1XOQV+yEJuIlR7dwqZnHI1y6vD1A2Q
5JParFpWtV7DTpw1/5d3ZAlo+MJOFQI9eRxCRQ2OFoMfS9uuywwyXAlUjO0GosYj
xbbv1bpVXUgPbXzsP6mXKU/hHAnUOpf1+osmVRjl+1gDFqckp9DkPWw41yfe6K7I
74fCU3Q/PavkspR8afTcpO6ERLl0Yfd5ZZuySs2bf9paEqlq637X6dGXmpmKNbNx
+fx9t2SaaaSrrFjU7oGPLPtSEduT8inRD/M1CPcU3xI/D2EXD1xBuiBx369H3UZs
TwuCfAtI6tYSyYJUFACYr7B6SjQYQQvnjWjLO0rzjznmZ4ON/cQNqN8CZeftDAE0
VdBdJy9P6GVLtcrmiu04COBkWbi3bU+AJ2iDzEDzx3J3MCUwyd/2Mr7mj26q1AfW
YqJj6p8UZKQ1QpTUvZbVg6CEBmcGp2fAKhvHHmVSQFAf+qMJ8ZntqPMnA04X9RLd
wXAv6/rA+xwj3ZxOwguFC2F8z1n8d9H2Ic/2Hp6zhnJ/ahY3fvr8fxK2TlPXx4BU
76Q9XB9rZd/LHKnSGDw7cSTEvplZu8n7cL+o9gijob1luzytZ4CWKlonUFSDJV9f
DN8uykhAiss+9++gC9UMCjcv8v2wygiEtg0ksENVN2dei8aqxNbmgPMMmqCc0DKK
nUMT7/TGnSEEdT+horBbH6KMWrCV6FEpidvBQjHULXcAbF6ZyMLQIruZRK4POPu6
jG8zgQfzlAINYunq954hp7dM6Zy2hGb1QCWJ+/So2ZeqaCGfoTkA9DcafKs6zYxc
lzslwk7G0bIP9gXr9k/iLWfzwDA3a6RFmsHVX5nIwhchlISs9eqaA10CfkEoWqK6
QeJgowkSSMa9/BCgCpRVFC2bSqlEO8SSruxT9oPr13loJ2mMXu9ncms0+0k1NUNc
53wg2NL6Me4Xq2RmP1m4/xLgw5N4aoMhEwOX0atRHii2kbA62DOZuILN5yKAbu9H
yG887qsRYfUaw4zJHy2BBPFrNOeI0JD4cqcXhWFrHyrt1IHt4Z/3VOE84sruBN8x
P9kSjFx7iollAXOwC40h0SivHJO94WLKir0U1+ZYDIUCAaxQJVLRjjStFbcU11Ia
Ig6xVcpW1wjM4Jrgh8g+hFdWGWPYs/yoODSEO0DJkhjyw8qXSxhOXIyrk6qlfO4w
4dVcI4pYwm6Tw/NgxH02syUJ+akQ8ObaT5ZRG09wm6zV+jQ3emAYfiRHxwS0nEWn
Vx+KbrahLjc2tojaFlz61ioSTfWeHQHe9K2i18vqtgpDKLlxbOxvovJZW2BX1Yw8
mrTcxqWMU2NQ/TBNiaqyxLlUKTdt8IcE+xIlySJ2qheWOuMYwImSsL32W6VA+DHR
0Fn1WyDX+y9MGP2OGDAzerGG3R+jSTh76xY1m80oKlRYp0Z8QtCXOTmY1iOpo74I
cnXqCyCyszcmaK79Ay/3hyMzIl27jVH8hW/ErGLa/IiB4q9blJTEQHJY/dj+pImz
HyeLxJOwZmq/qGBGQJa1YMHYEv/tQOxEfpYD9UpOmnjj85aILFSizAeP/xSmYXVk
2bwJBJ1vhE2r9DYsdcScDl1D/x8FduSJyCIkDzXVarFa0b4bK+HMWMkL+W7PqBaU
YvgcYcj3GxaBJd8xkjlOnQJzdyTtJGojsGaHs2bzBVkZvxwH3Mt1X9bjrEZvcy/U
kOuNGmurAIYUrwalQMSnl9WbLw6F5j4zE8AvXlupGRGZRNHjLlzTNLfCon+5tGhd
irnTzxFsGGgpWY5dLqD1R1lRfxoIOluEjVCh5ZPolLDjPmHdegggUAcLdlHgFC9J
CEOVq2vTcyyFiIC0VBO8o2xI6BS89y7IsCOHHFAryyOyXP2mwY8jACXxM/8D1Jod
1EYzkM43alZzLMjsfTIfXGgOv1O/zDGwZTMlAldCyd0FYS5M/Ox0H+rYftjgzt/7
ZWX9qtLPxlarhbS3BFGqEpSJQ6O/lQw56lmOzXoDjsQijGawxNJCILd2/B+reCAu
HUbE9ow1RO2e2+Mfj4k8iMY7M9mozG2XfPyMiv1t/lTgSJ0H5vExQcqCM0WXqe62
ZDsVnw7SXJ6lYSKywyTk8tT/l+WtM9l5as/Pm8KeP/Qfk8Gxrq0n89fyptEqDLVv
jt61OHPG/kx++GCOHXKWEPFevwxrNV/uiVjnZV9yxPaXqIxUF0/RnLfWELDmewWE
Uta4zJfxb+c92kRLvqyBqj6VpkIkiD41fuOmFpYcy+Zu5/4jmk/08GUvgdA56nac
gDQOKSHWsraGTlAMC6BUyMWDiAnWgqHPK5jYMbFagGLiFPvjvi9xGV+zQIdPYZUx
qeCTPgQbifb0RNuXt7rh792Pam3grI2EJDKU4QNUIsKj7ohb7CzbKJ3zXuWgFPJ6
nO0lc5v53CKnDZTs71/xulx3UNdFwHVE8fGvXnbS2Zme7xTJL3aP97h+MLPweVLI
h5K+joLmqujNrXwElwIZIAunZntmK6Zs3p/PIQD24wJr/O1YmqSg08nWAJEjiWfY
k0WgRl9RbTjI2l1xCluloywAZfbIUpBSYWHDAHxIrzDWkyr/sDHl2TYbYLD8lRkH
VM50VN1IBClBpyPNLvcGT1+wF1ODWviqUNXAYj29pzzmXyW7ljC+mMLlJxT/kILN
0EX00gwLWK3FcJ90D1YMZbS1aeEuKYOnRYmN9kERWo9l6vzHjcsmMe8+/wnfNtlb
MFHHlZWEvP6Qu0RgY8FNWA1w+M6I5wMo/jHvL8m/aUbgWuPzacky5XezfEoIF4HH
oS7WcomcmBFikEk7AwCvy8CASMR7ECOGbOeLPcl7o8tM2VINukZDqWQb6E9lUYg0
kSYrgQArs+aYHtxNdb4EpQKCcOjzRcixZ9sfaXT2t6nNffrF/CpNpj9uE+DtMssm
VlT63pexlLxFk63tFYfkIlZMDFlQ21Sa7QvqUvTT2nZSKys7AQXthRpf9rrcVGw4
dHZ/yw3FjvXhY3tMpap1C7SiB+0bFuENSo8eR9kgPF4pdFnXCPZolweoFI2o8K1n
REb+HeXM8erJHs6IA0I3kO/+gBeGEXI/P/IGqQjmcVYyrFBnSZHRZ9v6gMjd9AdL
LcRco1W1I6IPKE763aBEohxaQ6JUr7FEzni2ffilPqpZFvW/IuwLdtjpg81YZ77F
tFBRyTeQOQqAUrJ82bY2pPWQgW/KzPNkWLx2Kf2NwUDmFB6rkHrJB+uSPqnhoi5Y
G11JNdB+I9xSs/46VE+uN6kO40jlbnE3rZFoJVpJN722a5Z4tYeE9bpQfgKePCvH
4af0TiL7LOpQEHbKDdSwZwWlzzL65FSLaYa6cKACbjd3kqX/X0S+lZx8tjH6dMga
sNgKLgDDxm0c6h0ZHwY4uSLxABnZtiUtK62JJMkrEbW0kuP+u+53kLEiS2fpeck5
aC75qc3c8vH17k9wwB2D9nahlxo1giXf+fwweoxTC+ylUkeiYqOodLEWKBv+sWGU
yBBVdQloYbxXfmHoej/qo4WZ/BVhllGo31GtUaiEyg6EjxE8EH8auJsn9GAeH9us
CF/qg0egWN6ZFSJp3eMcRb20+b8Vbro6lMEAyhz0aZDj/rUbHw4GMC6k2EMuUH1j
qMR6PyEOsLOTxNXmMXxEChXXL0nHlQb4SVdQ/2V/QzCa+E6NynJUSW4OzATYq6ZS
SLeuQVKGbLqrc9Sny10X+8gmTJ8p+kJ5vXs+HfAx60vCgUx7tyOzLAp3WuRXs2qK
Z/Q9gFfb2VbO42bk9mrVaJZLx/bA9ZOGI+8KfFfgLThH8/qz+w4y6EdFZ2tKSCv2
SmEXetzNVFvc47sM7+wfhKWEa/SuRvn9Qw+/AlajVUD39+H5024DfSiH9j1QU6F+
n4THABB1w3ec2C605h8c8pH/ddtOIoGf5xtq+N601r1ZS2fiTjHoO2GKal/64Xlh
2A1hdyuPwVCUuPPTW6iGMn13AfTdgLzvz3ubrPYG/xScXF8cuqXN2KRHmFrehdMj
LjtlxnIGtiD38ENOnUmuDwuojnSX2FQzna34oAGdj2QkXz9D0ubeAARqFDBceqKJ
P3Fbtkjj0wggt1nyI2H3FvAkZPXoKyjhjJScjTBNjAjkGdCH7rR7PI1PR3DDzvk2
9dmnVy7zyRes+VQ1TbbBC2S9/sivV3hqiGNha3fs1dByYnEqWnGgDFV3NdM/MFFN
GbWiisn9Jmxi6x7WjxwL0D2V6kScvJVp+1g77QW2csD+Kk6Iru7PNZCVlo5chLko
VT4Vfriwn7ygNbcBBql8tDDmn16nvCkpPMS4x6XVGMCBWf2zRwutlyb0u7Sx2I21
v2lCaXAYY94bzRvhHFbwIPCnG0tYlW2gDwtBfOoYnnxyeUf9zmyASdQ9FBZvAqlU
4EboZlTwmVTrvp5Y7LSYmkQognQI6otUS+LHLwua+hcWvJbTQu6evKCrQNBZidJd
d+JWWkIhMNTeAPfgQChdLlkHhNGpiTdgVdnb5xNKaDUNTSxbvy86Ni+zJXIb21A8
pZ+uDYtrRST6evU+gHkV79StQX9mwvQPRQutvtg5aI5tDjw8vxjVdXY6XMMBrkJf
Zfq4AoVFBOK/zRa7D0RXuNyp8a59L2D+SaFPWIztAjBk/nwrbcOCiOdXQ5blKKpl
EMrEiy+jcrjtZqPa9L2L/4z0mA4a08QCeK1zgIqd8ZxcUCwwEROUS6CY/CZlyY1A
Vz7dNgl4MGVGBqc9eE9jVI77sbWwYW2o6gNzO1fnNAnaBDVm31Wbi1XBeCwI92MU
MeefkmA9LQAjvFBt+8tNQ92Bv4HlGO+XkekalM1HvmLrIC3o+01vy72ZLYHPLqPK
Mp8hdYW9NsBuRslhmETMME5xnlkDqW7vUNgZmTQzBBjMN7K+s3PpAu5oIRhMuShL
BUaw5UcqFhCcOU1vavFZGHX+OWhS3zZjhaIEbS51yy8Sgz/0SNJtzo9jq8Flsrlq
UcrWI4K7ER1vu3Zogw6iSF1SIz73cQznsRQo8ruemvZ/ymL+p885Ijq+mEFN2E8f
AwHdBkiVVV/QY2WlRoScivXqdq+VcYWqLZTd1F7ziqcZDdnI2u82xelBabKQ9/14
5VzfNbVQDoVwazqJLeSrW8pqeMaJoMUquTKBooS3YR3ScPQe4L0o/4j+0iBgqKeQ
riYZPwfwGrgNThoNGi8QnCChiE++rwm23aOwWqeVqh43jgPbYaPM5Nu4v/fjtO1i
4NMAE4yYflUdboesiDTag2D18pPLLTao/kp6XN5gvDU9yOWdIJDYSwz1gBAUbf/n
2PIlcquIO9sUlUwoMXOfnKiqZf3M8s2W4ErxNWOKBo5G7mNCmZsni1Gi03zDor6W
8HeOvtx/6ExO7gVh8nO65fxYt2QbihfkMc79QOJ6L43xpU0ngBLLLBsJ9wmhL15z
6DG4uQ6nPPjAPvD3NK9nZvaa2piRZ9O6MwuMuAVTJS6LO358sORGpgt+3Y4IGfbC
7LP9yn2L0tKOu56DzHFQbtCdGFz86osQ3Q+Um2M/uu7cPqJjsatNj1OEH1FEISh9
TojVjvnHLJFb+JHjqpd6dYsKdQvxsVxe+Qb3+uqbE+P0KAENpCPWUaEccpBcYtvV
7iH4zP+iHHjxxAOSSUZ5ETk+jLiVzCeVYd6k/lWsGkyiazejffTiorvrZTg646Wl
tH7xSO1acV6WM5qsNBx5SYmVMU/NRH9JUZMOB2TJNVqUcFBS3RBt5unFAFlkPNqw
EmAGnRCrZ5uChUpJpbMucMOr/n7XjpjG+H2vglCqyBlA0G3OXPi9MKtQT+nm8T6A
KGYuDYyKwyhfBuAHe2tQ5yN8goetrHdyb8jSM8ym8sgtyaAKSyq75xrTg7ZRmhey
mZOxJjmbR7svStdDp8H15ze75IopLqCYe8pfGeni8Eqb6ilBoTQFiQDpRHrYlSnt
q7jiWwLS0maca2dBhauOZau/JXtEniq6l40epQpRNB+OtwyB3eojLoJ+sGdULvpF
2HJfRjNYBPRYGQN/FvY4i2Rsc1Am55TJOAl6j6W3RqfA+rPt0xdWtf0nmZTcCghS
25TOw3IToatfTleCXBpIOKpEQvEC+LkV3fusl7EhAHaEJduLqokdDvaXSZpWHQN4
/u3Cf3zP76AIOJEgEeRRwUABcrGIVEfRoHeIf6+SQNX2hTYY8zAkMSQeazPwfSka
ypamOa4Bo2O8y2Jqrm6jLPKDnkmIMD5dXgy4wQTM7iqJ5rZuec9btd20R0dmtRqN
+J1+EHaCHrGVFK6m+7z0c2nN9ndM2acizs+sPxWkq9zgA4OIEwg5IqPMLVIA5EVX
Rp+7eI93U5OlmRgTl9HyLVgc3bUGRwKPIRio51PgcHtvkNCaD7ip5ltwTuYEEsRR
ESGg0c3bx9ZodlMUjcBftMNoLYHBBnS7XY8esjvesmqWli7qQea3QcFkcwVQbPfc
aly0Q3LSEQJ0YwYHypCJFg1b5nudU0XrTvtmflWwmEYcQ7d6dYZ81v0DwfV34Xfn
KTsV5LugTSlXEqi6e+ovMq5HVL/fHsmxN7pGW0f2WPX75lVT2RDAk6BK0Jx8VDfI
xiwyWu6bloPDYdaiTPtMlkBQzVLzYKkVcvp/rC046/ClwDa94pj5ZtkQvZ9Yx0Vp
pN6ya52jHl0+WclQKlORAMDVkT9img+yvIaPUr0MNmuuGZ10KANOxMMvl5KYMb7w
yWrwaTxhdWsLYa0ZEemuw9TTURvuGEMhCymuUJcJtf20VZseln+QK9nW6w+qENy7
gXO7HIJ/rZFj9DKtbOhG5Tt7FgzfCb9wXIVbjo8VLeKAMF7x8MhYs23hmRa9q5jZ
5NSyTgkp4vBJhQk0xeYygCXVRedf00cyv1brnwOynYzLqLylY2KOsPutPMRjbCJw
11BS2chKgtI/59du56suw/dzXDDYMpcc0c9X5xPWfIfzb4tBBlXUhv1Zrm5U1LFO
6ZB4kJtt0hShJJwSgq5kvciAf7ZizCSIlMSzS9trhw2EekeQfaI4qeOa+bPQiqjx
t+8l+8plsFAUfuUgC4GB3LNjSHP2SaUFhbYeH35aRqmrnetYfGvJTObhtNY+pRqY
woDO1MWzmOBEHmhSJj2IY8DvPxiwbyRmtDFJA5ZSmNR+7TZz2UigbGbuVtEqYSIC
DhT8OtOYUyWtsTCPiI4BBKkJJktxM1NYbbW5PgXhNkmTYfBZfgizHgmtgrf7MEDF
qf/rJinYdKHpst+m8jDz89vrGcOgFprAjfuaK/oLrMjkBs2qcHz0/KMUeeAB4v5c
o/jup8Gfe24OY1Taw3hzBB5hjxrV7Z4jgyOi8MOV7eXX8WvIs99FGML/W8n6ynbn
mZSi5KG2cMx9HQwuz5WV8Uv6/mktyqDXAxYco64nSVFnbJe+CDHKpkpXHAVx3T+U
d/VszC53MwsMwgpRAO2fJ0H00glWRkcpZhrMAEgArV8U8ywN0dCs14+QQNsO9bwj
zcN9t6AwL+7DYNjj6J7RipwmBBXy8hhtUGUSHowrZHnPCoWsCn4DCiyyJ9ls4AJv
nKDVYqfnglYe82xJgq7kkJoPRj1wijT2M55YanoIXgX2Dj2zBfmd1Sqso5qQsSJ7
p31SHL/G88PaXscNy+BQW/p/EWI6zvOrUQSUxsxGHBSkHTD1BjhqVeSK+K36UB0K
wf8inZGdLEDAPuRAgoaTPDpt9cTdYzamGJpYEa4HeXOOJcZhpnsjORk5lJULQOKz
eE0lx9ULe6F3OzMJYUsRXBesJSDlXHiC9c5U29lGsZiSXAGfEhqj/At89Cdvv+4N
fF6x/5GXsp75SfOMPbd/ozff/Z76pN/hmqvVOaTc2xDcDmmdRlMT97F/88N521FJ
PhDuBsaJr0M5Niwbh5ospt+lE/ha7IwsEpOUsRkY5P4Ps4WkzglyvKZg+6WjF045
CM3+djbMewrSIqyVCAkmdtL4pafaNothE3dueUpmzXuwLTGdKI2GPq+YLABeKxUK
vfOntnJp5S7UZ04Hx1754P3Ewq/CMQJM7u96UwT9f7iiFl7csJyBoHwLbnb9WYfb
vxi3x/pDvvfYcScYbcqfeLpeOsuqaK9TDsvr0L6D8WdAaxF6vXz7ugOBPFFPvNZ7
5ooa51+VcT7H/FqFZS4IdWom6yyHkweC7U4d4QmygGXnsNx3RoVo+kTMNln4oKxi
fe1tEfsoWu2VaGw5CLxeNwXCw0Ik+WqHTZgw4BuJZwZ99/1Ni/BbaOsEBUkXgfWD
103JcKSB4XQ5lRT9nPlvZb98RBZKMM3A2L5kWu/739JPjEIrWcYKiGddFonLgXo1
iG6katX7DSPFLyXVSRBY4LA1iPeAtU2SqV8JITZKfszPzEPubA6SkU4cJXbVQiwP
c3/5fXWnywPub5b/4lYImf+oPPK+B4InW8kIcXmGMWUAJSOfMQV8uKxyTojgb7fg
oItPJe4t0jYWFl/R1sZlyo0yppoE7QGSLLCnv/K/yYMAR4ZsjRF1GbI30AfLthsl
27xf4b9HtCBONA15qi4qDM7PUWMFW8fIRX6eOeERvnkXW97d6rhZZ6NQ+7Cxk8iK
55BXfRQKUkKxuGge3sR++xrSce7OQjeOWeayTitH5gLlUJ+GmNyIA3NXOh3AbhZ5
c2jgYQGSwPDb/XIS+TMiyjmgi42ax6ToF/peyLi7/E66e6+vuB8oN8ag1W57mat6
Ny1FkPgt4VhyJi4VyAyN5z9D7q91bCL802hl/c1sKPwQuVOTThi8oYDsBD2nxaPW
ReNRMzuHMQrgdX6aZCWfXA3KGTZLDq02Q3okAUK4VIRT25rPw7xizhXIy1UFKY4T
csGAROsoV8Xz5BAEjda5eVVnvw/Ac4H9ZD8aI4/jSpdLtBE9rINJDvBKYqsW6aLd
0nr/YvnI5eeDeIaZIH+5bAybZVYqK7jEMu6LtoHAewxoV0PDywQQdyN2du7LhyPZ
HBUOfoM7vA8tgCsqjttiLI+LvtjnZCh2vgGLcwzhKgF+vnzRuwsoj05XFl8CN21u
PA4yN7d9ygu3oPuCu/keUGBkbA/A/WSTRnFUr5RxOae7470ZZgNqu4KtuWPzUurV
OzuS8M7SIXX0qEb/YVIjqI/w2lvv7OTIqG/gamTWS69KjGKCjduFgSM/VXwZPmMn
KcJUGHT+Cb2aRzTH4WmtRre3YNGSHSk9C0QLzJ6WadzbvAQW8Y4/2pwdWFjye+Bg
qvWOHc7wvH8JFqhHjJMUSENb4BPBsTCrUywRxnxv9SQZLbpNmWYUXE18F8U1Ln2y
pco9BZwfdVPg8ezqxvMTKuARaD21KhfkeEAKBlhwPVze1rI5sO5xBVqqwkB26zBC
mzwqLUZGYPII8/IFBc3ESKgUzTXZ/xi4ExwF595e9pQoEbFp0o1Gsl96F1vQgG71
BVxi+aROSIee994i81fe9DL6lazWeM7vbTkfYMkcg7Pg8NvWpTb5jbIXlHUbgcVR
FOYoC0hnim+xzjX7yUGqXlW/++r6AWwJ590KjVmwTpfM5vKPE3JnqQ7HqtA1IBGJ
0ppbPGV2nuKKWuqLz0owcWohzyKOMF6gy6tmxxorgAl2vM9bbFyjKU3Nb2PqCmv6
HT+GFUSmaHWlfh7LRg2/MyDQABszk5p4IDYiO1GaVwUO9DT8J6P5ugfc4O96x6IR
TKPsZPucsNHWfFMqGXFNyzL34cqSyhv0cI4GJ8fjk2OvhAWoYZvjQklK7TW5KBFu
mmGMFVR6rPVNdir87TbMN8fvjnobzjI54dprcPSBt8A2FomsKVa1wkJ3R8s2W35C
sWVSiekIKKYckJzGcrIyBJmmtD5OPs4PWlSIulvpJwMvXhzD/udeeJmT/Gk0GEaS
T4FLQ5C+vJ1lLwO9CTfP7gtL+VL7GcYiCN/kXROfxf4Y6GdWJqmqmbIVjt351Dy/
ctziyQ8VTkXe/mDPf6iSsZscMNOZLS7BGvod4wHCz0wN4r+VH2Uk4ujDBiVvjp7c
cbqg2bxLMIyKD3pWYsiwn1/2+RXDLM6JZcDNFxa78GvF8SYaVDCj/RQ0272Wg3Wh
baA6psp8pNihpzOyD/QtI7Mtf2ETKBdWa6EWhNDWzrWfkbCvBwoSda9QJDyyAJ/4
LRsAvrVrOlsWBrbKk1kmcgEN65Qh5p7DrZAa2Q7NA22JgKJkiohcbJKJmtfvQKXN
P0FlCZxwLX3B5nQLyalYudgsZ9A7qYWE/2ZoF1n+CMvXDi8VWEEFVT9NkpJFQ4eQ
LM9dA9bxmDC6pr8XZ7pE/QfCL58tqsw3m3dsqXcqVntfQoS3Nk8lA9eyuYSlhs+m
eYh56ROlWeuMe1xtGJN2lay2lxvjlYyqS3V+nO/n+4PVKHeJSG+YqYoJXqbEQD3t
eJxMXGdE+jV/MtMvWmATC6NFMCB7ECENOuvQfvII35cakFeMD/PVEOvumpbUotu1
m2+30Pctjopv1lB52pBeVXJSo9cgj195/WNIVHvaLVvrP4zDZKSz3SxkclAK9cfA
XCcJMLehJFWxIiR4l/mJCMOpyfw3FyHehp3KY7JyifopsUFYaOUJa4FlOdmNoWzb
r2lPw6tZ2xxSqS/OttVfokQ09mNjWdI3fKKOfRUYKmE+ysBBS4hm96u27AB7rAg0
DCkcabBQavAMpIB3A0AzZgLOIybz1WglnRyjKME/0BUZm0YR4EX0KtSMPbgXBMap
rI3bQ8BAHNN15oFfuqhDR/g1LwwVBD4+xOWD158WiDTXN6xH9JYcasWpyDG59/Xi
uaUPMJb6d7z0xOZWwVMSePQiqFgaKoopDcAOKJkLtPy2GZvEgv0vlHeEpTaeZmA/
kXadPQbIZvR7C+/3D39NNe+p5yDbIZoG4QE03/iaHsQCcui9/2wcnqBwNXR8GPT/
07U5AjkA+FcokfBV6bwMPAAU0/XGQ7Zk4WXkE0SZmLtpyM6zkFOL3Kiis0gVQInF
nOMT3ayXeEtpD9PABy9mIbs4Ld4jeouS/FSj1QV2q2WqG8hv/Uqq0TwwZYsR39Gl
GGRMMvVl1H8dCy2m0wGD53VdVkylMs7LhPdwUl6U3cndUgArbyeBzbs0aZIcLNvm
5r07g4K9t6/cfrlqq39u8a+NnsvfHcUvDu9xziN+XMKLaUrm4TGfE9C0y3PTrhgW
Vlw+dmTUb+m3XRz9BJz8lvDNO3cWuC5DNGUUTiIxQxyBnG59nOLVblB/yNQ8KYtf
FcsPvPoXkg81Daz8r1bbQ6wUvCEdtS53VZFQQMB/9IpLXo8ORb1dE1s4IA6jX0tA
3g7Y3mHKGy37Mkk6/KPxwqW80m4wk4dz0ot3J7thvnptW58KC/tExHQ5/wlRuRNX
FS++viFr+4riE8Y8cXluRUdC/x4eNX3lI4ZdtvzerbKiw59v2AUU3Py0gAREg0un
1XJUST39955Y+5xHlgRCJNMXOe9hIbu2mi9x7FaKHRa4a8uyKnUoSEbtT3RLcRhU
bjWC9Jfs5dP5jdRapEEU/RcoZsHA2ePFaitKU+7Kx/GWc9KcFXUchW3/6SV9cbwX
8EPo6o2+u708QDpt0u5B0LU0oLPqcz/CO0oZKg6kvjjmJl7iodW0ynYHRDJtG64x
bChY9zDLIVQb96dHJGu9sHvGOlaYIR3vHvIgztRS7f6KmlMgCGFaBI4flPFDP6KT
VFYUhUjIUnKxb9nZ0AX7emuIn6lWmo0fAANDRy9D1x4f1kMULWajHMz3b7wLK6Uu
TrDEOqjRoNgNF4DwpyzerZU0n4Rco0mS7rNEHS89vuyNoG67etyUE6T00hsrE1H0
JQnFHsbbdQzj4RMDR9QkItV+nrZ10C84PXZpZtvqB5UqQrxEX0k6UsXOkIaMLZ35
pmVt1//iZWUUfdOH/Z9dceH1r2cgLCNXxKUyNtYizDjiydCLRA7tNnSIYXxxGj5H
PTNsnBZPF0Tg8K3gUc2K3ihgqp4MyW5luJxJ6nLhcZivweCy1PWaG8zq8gxt+eDv
we6d4JniYGaSU3/RsQM2FHKKKiCqEQj6/KEEWwS0oyY6lK1Yp1ZjGAiPxdcGf9Me
RnrNElwEG3mvz411crA10ceYzWYsXk9+oL3RYH9Ax07AFdPxgWTzNir9sRxB5FKo
B4iZ1cn142RbxKnH9flCwhAE1RDVGr0npFlM/xShf0DUYgfiG3Nju7fkkiY7yGBK
iwHODghYp1d6iNAwFf0b0nEHIsizrmonwCCghd4zXM63yvQkV30oSbNtQQlvrhTs
Km2W4PCURtHDP4cl5tdgJKyPe2mrVmNq3PdHHqVNphTx7slYA9ZSbboyQsxUcahd
3g62tbnpRAhjshpY7c9byb0q9126/g2G5TrWYKwnlDvD2ONObm0/7f7MTHfgYIYe
5wIKNKSQCxsWXWPGgvqUHcURmtvM1PBjP0XV3YjLtwAR7Wqq1U90Rs4BRHy+ggLK
eRGGIxvkGjOsfv8fyw2Cd8yb2qBoSmpbBhj5GZjvTa7j09zK2LDEZKn+RwAZEGGK
z8pYtty3jDB5M71mr+V6fgwm+3Cdc1E9NFu/SVktRIRHhG6LPdhZqJLXUanJk3/D
O+v4ZfMt5sS0Dr3aPTLxSzAfCd7Rcp3b3XJdTTwKmaFBrnkKlL8yAP6Tn+ISGXRp
sF7aKMdsWYylUeM4EEaBqwhDC/nHKlGoff1f+yr7RSzTFcqC+YcsqHgRpQAZCHx3
QHz5gmMW6eC3shqwafhuqAXd576hcdYL70SwQb8vM22J7SC6jQF2OntBDfdSSO+Q
VZ4U7jNouQIrxYPfvVglAbEnvDH4Y4hb/cdI58XqgGTw4euHzV+/8mUcullyE+0F
me2fEIUO+cGdCax//KVtJ4sMSDFiuJ5i2Atapy/6MCxvn2WNhJydCL2kKXbdBL8f
KKApAyKirroVFnvbpyou3Zj3/LGjrXdYu7ZViTHRG65rluIIPVn+4GbkZ5nd+6wP
Ru/DYn+EaWN/o8vEud4xmqp+s4aTaPPrW3BSMkxJ/s7CZNZJiqbnkfBY5j/xymAE
Ksc0yCLB0KlQKax2EwXMVzrIa2df3HaHlGL9y8KSahRXZ1rpBagaBWEMxcGduBGz
u1V020EEFtKbptFH8WOYEr7dxOStHJ92juXlCAD+dP1bjyOAMqz1YInI4wKVOt/3
e8gWgR5iSDwV77hdNDgN9lXDAxXlSy1L1QnhxkhcVePbK2gvGNCdbilPurAj4kzT
mu3rfPPzEA/YDX7lGeYyoRUbnCYMan+F+DQeQN8KZkZpBSLyTaQpHrLgLxJzagnk
ZnK/ztAPi6DooBg5x3crCv/LuLd8BpRQKOW9hrtS3CzOVH0kGLBQ3AjTDD90TUjO
Di9loogzYI9YcdpDsrPgM9Jlk+xKlJiyZ8GyGnLd1L68pUme8h0ph1fYWVt6x7mc
b9gPkPZS4WoVG/lxcSLCdg3crNXg0XnrjioDe8XBhe7iFEKqcvcsmyvFJ5Z28ZzI
jy0Vs9A06btDHkhqyRqQnmDp0IHaEqLP7RpzCnaGhJQ7ZYT5LomZUUSoHOGiMJzT
DMnjfcWwoxYnHMtb+9+QFF0MiojcSKotY0Ouxh0ETM4JxLqXynX9lBpQ1r4mZNyp
UkympATQ+kodXcdPFd5E/Flhmz7VvepPolLil6ZS81mMZ7l1Ela2QaG8Mbegs9AD
dz7Ijh3iEMHwCb1CwX4BouSmM/eVTFIdX3EZd4MMrJBz99JLekl2WwoNF+lB+NBb
xiDvDfuDhGduu9nrYG3IEnGvaRpY8UeRFOGSlN7PG8HvdaITp2zYTOWra20njDU0
Zf6HZiL1aVhl+Si45vXgasGxdeKCgehZ48y9FncmnvOWR4zKFjtdE2BTBobfbiAX
nBSLsNM6XQNrXfLdqf0RsVt5PjgQzP2KPURRb/yskUop0yXQ7VHsvzDyU7axdeRW
GWtSyHPVqr2IRX/qimUBSNF35IpCXv3BL6G4F7ABORD7HY4Ki1j7k7T6hmWFj2Nm
4lmu+cU7KFBHBseiaDPBG2c2/BQ/UozbAT1rvkVM0T7KhH0oFeTBxJmMSoynXUjp
1yMXJAFZTkOPqrCNjSK1lJHIV8xaUrRxfDYWonFrIHZq78K/pYg/+OHo5YYfYTfk
xiZeerKg8t9UweD1w8ZAJMFA8XcUYQkL/SOdyVnAuelR8PELFROEk33alDS1H11e
YDmKyjKHmaBpAy2cxR13e6N7/X6uXGQvFumKnlVWWjlc1JKQ9SzEAa285KGgq6gl
Wvg5kg4ZU4ROmqK0mq5S8pCYVs0zchyMleYKg9xhVIo1nosVPwuH+4ZrwXFcTDef
zn64bI2rQkTmUcdjSz6/2Y6RkfcT6U7paQgnM2d6uOT6cMh4hY07Vy1tWbH2Qkgx
R64ajVMsgmrdR9lwDS5iyVw2XF6iSd4ofcEb2bXfHY+fjbTZ1PxlSsT1FzaLowz8
ltBaMMt1IgclFz0XGxRlflQmm+Sq+u6W46iX9GGPzNOXi1kp+7Go1URvBmP1pr+u
BK2TNQQbCM+owDJXhvDxAKSdBCUoFN6gF05KqXV+Eo4eFWvnQW6pHmvyDa63o/L/
dfR8QplF1apGf2AxikYTGpazd/8eLy0yL6VFcYH/gkEbcD8hYmqcSp0xz3rq/rJ5
8aW0/rPHuZMWqPu8Pq/vLdmrycjcltNUhY5EemSBxrHBwl9pKnccnx+GQdODQm4A
DBa66GT/m1uOZG0vuZTsirgfzPHRM+U8b+iFh2LgcjgVC2jOWQR0wR3E7rWRZjHG
m9hEk2Kzt8I9+9r1yjMfsRd++Q/Lr0815fSSrQq+6nPjVn67ynaUgGDsiWZOKJZF
+Xt6ShFLPud9t+dW8OWaaagdiynIzO4OFc94ALUrgMhf6y/BASCZB/oL3QoGYbEv
R2fZp9mlOVRObKccyc/YOmGdRpwpM1lBigjnGfuLqHxIftLD+BdpfYTMoCqjitOW
1Me0RDYA7TGqCBEilvoiukNcE7Uc4U7lI39rDzldni/fJ019xkfJfcXhe8N+6uaX
74Fprw4n7ZcNn2ulLHZYR2yXCMonCHOIX+O8m1aPK2mAAGFbsYt1vOrlyKhFcFIw
swji9qFWP4xQeCLLJ62HN4fiLhYLQDj69O0KdFGldf3ilrt5wDfJIKO59Y9wtHMS
t16oYpSF0FNSDqsAcs/DcNeEsx13+8Emtg3Fp2JKMqFfo2ZEXjchMcn81taN/RcN
yTk1SbErw77keVLzNcsNYCZTc3V5nNZazZ6EW5IMC8YRSru4lXYUPdVz/FRKlZX2
r/dtFSkQoE49uvnJPHXxlA1Ins/MiLVyDehSLYOPPR86EzGOyFire1zENoCDnG2+
N3XDE7vEfeAbwn1vVWJ3K+HLPvj1LT1/tB2Ph+fXFlYakhaTe9KySnNa4j3oBDsZ
5VVTmDbQrLRsDsTXqJjArG3iAAwIsy+0hdfsYHO9ZYuGyJbDhHbZaWJNaAsW6XfK
2Rss/MqCYXQLA89hjsmQb76hSPQy1/r2NtWzcRa0VmkLVW8iPlpGuGSMR9a7VT2s
Q53JBtPvZrlmI1kuAV/wapNyCXvTqJ7f7L3w6ZKFU7ISiij04E7eRDkSQSTlLRrC
2ym3B4NQPnXAwZn/3r2g53bs281Ug0xGOG2Bv1jn47Fr+GeDHwF3VnX1AM7He/MR
LjgT39Tp8nO5yUcWF7rmGvvxXNdF7CQFPIZH7l6m9nxy68tqTpOTmHa4ZS8w8lrv
NC3m0U+HcHFPp2JGPwWO4nYGa/sAroyYp6tzWmnRiig3q26vGCFOD3pPGzsjlUsa
oX/2jx2CoU3lppiwZxYP8Iwdpk987GIe0P06hZX0mabX+4yQbWHWclhVrJVGk0Sd
Rt1qH4YSM8iRxJD07x4JuKQyVonLevgppxAp7vETrLzGDSNHSNQ8+fWPpUamR2xH
HFWTxDUddu24wHibtQBo6dqHtWibis75jy4TK+JCyW13XMzlTi3AFHv03ELc+n0D
DbO7dZM6zzNnQ0DYrkOy0QmedgAk/AgDWKzKA+cS2lxzXyCUfLS0+BfJWc1gUGas
IHyydLXcAJSfGuaVUGNdQGsDWoWzZaVY39TD5FzkmaEtiFPkOtf9WrYstgEaCx02
RzTfOBaI6mW2L9f0cWB53CB0yTyKR2iyQrHHd5IZ+ItyYxRQxshj5h3eWKw9hpnZ
ETsCUQH7zCqtq3OPKZQMBDkpyFx/H9FucQdP1TpKSDc=
`pragma protect end_protected
