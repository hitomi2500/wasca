// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
E84ZfJP0bhkIJmmXidTnQHqQZT4IeAZNknvQU4QOr8ihea/72YgBrkzCbZsEz53XDx/HESdGD9va
KRe6o9hf923FsvTx93N0rWmciywJYFZd8Wl07wMqAiUvNHZE+4pR6ykhUcnCNTMRPv/tjJWnkfns
7gETa9MOTX5tfEAfUU8pFzVPjxjty+XhdwEPawtASMwci0WE4gKzwgWotpv0Nx6Fe68lPX7Sd/hr
y2ALEP5utKvVGTTNZ3yvzoIf9H9MZlCb2GVaaMqCaeuvOzNzJnuTFA4DFSgfoMYum8zp6xyuPYgN
+8K5vrb4IBctMxWVTJP8mUV8uVNWI6Gc70o6cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
iJYKLmmRwLALwPlCgvejWvJ5CmyvqqWHMb+1JAVMR0Inq3VuRedbFgjgpTjAKIQ5+wtN7LAgjEJm
/kuHGBFhsuuhcSKWFR2IOVFQ7bo7heFpP2M10SajVAQNTDU1bjFUA0X/7rRwGO3/IUh1c9ayTEcq
ehdXoSNPv4Oin1wQvXnSoh20QECC25RFM9DUsl4Z6PxTqrAe6MagJKTj4+1u4jX53ZBM0pclrtiI
qt/zGyU23Zx3BKiw7nhLVFtO0NGdwIjXwdYhIvZwvUZhE9Oj7/LuOBgMzenIwGns/lwAAz1eAROv
GKdNUVT76QFAHh1cDHQKXV1JHFUDSisGWRhbfs74SuuvrwoB9pcxOg+UtC2/Rj/as2/ImvDsTcpA
ba4WJ7qTlqZtNIOeQo2ZzUVDh9C816LGGVVxUHKtdG1mcaJQto7OEVO5mdw5cUwLGejKWwrBorXR
6aCQfWd6uGz55bW07bbf8HjqWifv7S1Dyh3rmv4H4zel1xgS0E/VYyFNaXKTNVgolQ0g5ODYIztt
kpiQtLiLT2EuZRY5P2rl+BmWBhJVsh6+iQHdndrzkXExFO4UsG60Q1YfElgRWUPJG0p16qTdO7+E
fBmAv+9I1lMMwfB/6hBUVue/k/1QlN8rE3T8MKMPOYsizpkyLvZXc8gi+mBchqyqXP9PCFh5u7s7
iVgstOm0WYzWhjyEMR43Wa5JxsBD0pEcHTZpOrknIinguasZ3ws5vnH6NpuXVYSkwggPkt9kRFFM
W6dFxXt/Ebv4W/FtbsDYvgPd/cy54PvpfD6v3ilc/o/PcnZr+IWSzbnw5QtI/KimZiaXHhe/58R6
3CHzTDiwIs7fZF0wR0rhV2lj06xh2jmFext5rzFHiWX9YBa6IBQgbBS0pVek/I7yRw0w0aVEh2H9
8M2DkZUYBQr7OaOx7yGw3E3QwZGXqkT2vogEDr4o9JgVjLQt8OyQxmmliU/9Rtw0m5ov1OZRW8O9
yv5t8ZS1OhX8jgItwLHMCtdgEwDCM69DDJSyS1KS3GVdv1UBby4yF5d3jKt1FTqHaPTI3o4/wUiw
VJg6JDzLB+j+/iBpaKqPP3CXIgEQDsZ7KaufhaeuRT1tt2BZOK3S8CnnUDNvjkwGTxVsRUEhOp9O
T7ObjJENSvddkxpMcALzNIdo7voz2WPjCQwAhwJDKxuv2Tw40qEchYOxZm8KaQ59Zdk3zmYPZLYK
UUb9jdasaPxzipiDdyP4PAXy2BE/3z6CAAxt5u8X5jvHV4kFY7d54cKcPQ8CyvuXMh0+600usJjl
Ok7qDj61uhFUaDCusjSs2ogM9cj1V1AC3aoTV9oYyIO9N5j3s7eNAJkqWuVNMbiY5vwgwSG4e1fo
PUckC7naNwdZ/yov2x0yMztPMo+FIKCWmaMCnqxYS5VCCFKJrwHUFjMdPI2DBvXDN8aImxj4LRiL
C437ihKHzLTxy6fMPBXC2yacVNOIrXLQxR0ijVxwsN7vAKf9aNgAce3H09B0azcEUkCBO7Xfe3us
B31b5FLGkk0AHwvgAetHLVOwy6WIHufD7r2nQKGQn7lb69efPBx8nn39dnGYadkDym2gw0ar+HMW
QsGdAF5rYDBQCyihIsstccRq7yp2EtXsN3PLysQlkPsGweIMl/zKqaJGzA1U+KQkHa5YN5wwGje8
ysMMRdpPLH2pC5+QnW3fOx0TqqbRSjPfXWOtlG9QBnbF4Tmd2SrG+xEph6jyBsPBIV1ClL6OhlXL
p8OJwTBN2NmfwyrfY+r0xgNVjyXKG6E/GZeDpbUxXwqucug1YkQ9V5r5JapUKH/gK6A6XALF89yg
Lfs2229vOifIEQ0aWF2HGWhxW7bNaOM4tgLBTWaVkulZ69Ly22f7k1UyfOquHWct6DhrReVS4O1t
TYg8jszjUNeFHEgyiK3s2AqUuvAnYpBWEQu1Nq1wnaV5wUPbTxxrGYm1T6J1KCmSIdZSpDcbb9w9
jZlt+Bqw74MiPBDJa1cDep9rHcYNKCZomXSwPw0/+SlkwhWJJ8sbRRPbcwiH3LokYtGZ/XaujVk1
AsiNqTWqHuY1sdV/ytSBOOJU4hJpxuRIDxC0RqI67v5sGlVK8cgNoQLtpw4jsuFM2Oi3OI9aTFBf
Z30OJsyPXLAnO3rBYIPx5R+ekmdfBF91cPGi7b6D9plZF7GP+VEBtO63ZcB7BBs/GgY9b4Ng2jXm
a9RkTr8pCQmueGdfmnrSO899fHjqy3BenAocMc8S851DJRJ03S4MzEJT8bm21vdtCWoQcg4g6tUJ
GsPd5b1i5TuijbvL2sX9JkVDp0PXn0U+K9Z6fIUWpEeLwEnmxaI6mGiN0P0E0jaxAa+Qnwkf8VzU
U/oMtJdjbjaXNlaCG/MH2iMDThFlxQw/H8c8aUj9PGufIu1tOgzGvFSdYtnq0ucijjITcvKzTuiJ
ICuOrocyDzdPolNIIb0r/6GfHwX/WKrngnfWIJ+px7fpFjUkWXzTOsMEtxcdJ8d4AFdA+aEO2nqn
8aB2ImxjiY1BYmmIqc9nZ2gOa6HGzdbiqJbG7pOvELa6dGwzApAx1U+E518wwmbb0hGPuolwyKVM
J+FimuMGzFO2sCZzkEMrniyjAnSXyLySgm7koy5ZkgNdADRm7tagDSFBxeHHwfHfbQ38UMPG9aOn
NldFGHJVrIrdMCuNGkmHRVSnXxnASo/HC45q0Q3WDicHuKuj2l0NsScgltCyA9i/nNC0XEanF8EK
hiwBtexDS83F/X1QlRg4jj8Nk8E3Knf6NwD2Wl3rcwJvwJYS7FcWmKzS9s2U266Y4p9bSquq38C9
QUlEDA0LLe0ohg+NSMZFBY7ktpKpie0yWaIOamn1F8qpvYioXqR41r+ttQ+vNrQI+ZbvKeWCpZvR
rxTCU6ly0UAX67Xq5EO35vdiuAD9Fq7y5bSRdGuY3FucjZLqR8pMevuGe9deH1wsbtDmej+D/5pc
zPnS5ZPx4b160y2eeC9b+WAbECeHLgI7SjwrlvKnv3Q+W9MT0d4K4Ee7nPDTVdPPCO7EKnuGyoxz
zIs3ADMJ9Xxx7J+snWDP7CIsfJEovoVyfgCcNmd1i+wdvPsLrIj9GtjA0UaXGDZ2Rvw8hI8HLVSX
SJgsR4eYeJ1czgZtb4hPz1mS7Z7xIk8VqLt4SfURhErW4xQNAEgxIsNXrg8gYjfkbFdvwnoJgeqw
Tayj/1+77R18IStGmgPqfCaBbXclYXxAlsxokjKCH8CRNEUxozk/MkBT7L+bk0nBNFeb5j96BtO8
ohWvlp6D4zEbLKhqbVdtMgPnuJGVQ/HryMY4NdgxGMLw8HVqZsuHEC8IIPN2R66fmIiKciDMjTab
eM6uovyuQSF+zUWMlohTXLRPqDwbpdIXt9mHXz+k6WLpZeyyOrckISkYmC5XQUOFL+keCH0Olyd/
8r3UETQHPmjNLQjOsU/lcot0uQe4rc/N4NHlHsHZTX1lYnQ7JxZS0OuwxC37FL/S1FR9T4c9yQaN
PZzRr1gW1EHWUUFOvMGfjI/Tev55M2Ivqo2Kdk3te0RChtSnmKHgyDwK6xQ6f1rDbuYnKRJk0oDY
4LJ0QVsSm0QRrkGLJUPt/+IiMm7io4jiD6X2LSEyBV17g+v3yxckFGHa4kinpguet8o8yF/RzVIS
q7oqHUeLEq0RS+JloyQtOKd1OaXHEY+sHdP0ANTU8QlXHWKe6Y6DtbR9qPQbLOVtZvwY6lHR6W1W
Mvnd9Y7ALtaEROvmwAypxRNqzSncWgyhhPWqkgdZy4DPLlR6hG82Db8VIJhmqRRhD9n0haPo5nrx
nbguE9ti/3BbZcM/xlKpUWOR+DTQU6nK0ANK63l/52quuB7EL/02AVpKwkeyQL7j0szxABil8DC/
SsEyVqmIZtRpujKhJ8wRjJne/SKm2zfw5d8EDCjhYxGnJkq52x3wn/uGaPY/9ww5ofpswwJoL2EX
FjCvTtwsNp/bnsCN6HNdLl+fw/MDk+bBdX6RenMuhFEzvzXu7Fxf0cKTYPOZ8vqWqwUMGvpL4ZZf
9s0pO4kBnw/9czwZS4NiOLaP+neqbXeNB8SD/JcjqGSffi2DSXmjEEqm4K/yiK6+7Y55Ug5BuDDl
loqYvKF9MugLp5Sza/Bx0WM38FIB9Ax2+LYdbQ8fcL/WBJrCNw2TvUVEoXh+DHATDxF32s5mBEeX
Xzzwbxj/pk7RgO0+oLlEYeh7jvYEA7RcSN4AzyL9X6fN8giYkPs19C7jyNNWA3DuT+WrR/+CRt61
8hIa9bmTFOka0LZ025BTnCN5kE6PV9eCUK2jOXJYkBmApN87OIUHjMra9g7DOqlYbPMHYZbLs9n2
oWftZAPdZcjR4O2jpIvaiyf2DgsHxOW8aT/pkU90W6kCcsb7Y8uJ0sMAHe8m5CsJ7Udk/GT6xx+a
7OKrQZB1WdLLxxpgKiATsjUe35PURSONNK0a/Stm1yvXZ3dfeKfFVdush1b14KFzGuQ8bp+rxpbN
sOLq48WDm1s4uVeJ9oAY9aa1ot6lkpLSSrVhtU1oadzt8HD+QDU7E6LRKXfLFgMfZ5LagnFVgj7u
7Ah48nXPpc0QLy3COTPJILYiwGkpQd+fX/hEc2aoPkMvaOgxydgpCZu3tIE3H50K3xiduugrluvw
X2RJ/OUWwzx8T3oSheq1hPRZhbc80BUF3bFkM2ZbhW+V3qcXtx1m1OXOjv7JkF7mcIBDcFd165ez
v4Q5e6xO2Ta6337IRHzMouUEixtMbZyOlOpkvCcTol9Qa1TkvnBSxzXNrVng1h5g2Oc3uIjlYpW0
EXFQgGrvzohl8Rh1Sya553LwyuhG4/vI7O37Gl5fN0gkud7ixGNxSVJb4Zq43FhOsf6AX+0DHmrJ
ND2VrZrheogsmN6RJSvM44myACyEV6Dvxq7nigVmkWDGwGDxY8/OgkK0kleHdAnI5Wz3DwraJo0y
pPK1nTQ6nskrmiBG7l2r7RQ+LVtSQqGk4NXoQ5V0RqIqHxhSRDhQoAnha0bDQHhiZHYQ3cBYI7yq
4RXoecRP6cmUXpnOke98QpaqGUeGu1pVG1+LU7ikL2/QQQWhqHgvDYPzpNXAebZYVqCEqiWWg4pa
4lohSFJCBdcizfAq2nyA5q+J389ZGtLCTXWepy2nyx76POwPhomyimND80szQKy4E4wAVAUFWxoy
37sPlu/Of/+0DpPFF7EY/cue6DBy4d8dcogTgssMlzDjTFsL/qoeiMjSqAXe08JIiz799WmvL+YJ
r8R3PfwajbimvB6Z8rH+92Dj/xL5K7I8DeeyVIFGJsRoFewmGMWqlbmjTFCXI/kd7QKuQmsnLQjF
IjKF2FwYPhTYKOefFybwNVLlq6KPo3LmbygF4Fb/ss96fzHJtkxc8QgbOWU3DIdJzZ3MQjFJw5CD
Y4ObCxiHeJ1+sAP+SRwhgYxDoVrlMTCVEpoubjYrcm95kzw2bYb2kd+T9Hda2Vy+9u1rSJMzDYQS
KvmJ4WmCsobojkF94QxguL3kaZl6fSVzBHUnKpY+DRNGR9Pg8S3djumedFrHRxlSIeB4LKe0+9/2
/qxychpsl5iiaZxagA/wh4x27BllDCVe+uvWCMEM64/DISUxaLC8/V2TMYR/3F1xB2QexjZPfr5C
TE/ENi2Rwu6NLyxve9LHDoxzCW1naZbQ6uLLknKIN98Yy8yh+tke6DYArMl2kbty/9LYfa1/FTKy
dfppc07RAt31KKrltyccUI9YBI7EGxsBWldDRK+ru5B2501Et/2n+XEV1WmFwxiCKkb7SSxQmx5Q
b9WAnWbbPeDZ2tf4D31UIBkgUA6Ruz3bDAGOSmOGLwzjsEUQkc2V1uSMJQQF253ETs57gnDlUvRV
RmbZK5vUw6naLjzo3S9AeXDCbe1+l0rghId1+fOir0aaAh6lA6HKpI/VV8g67FIgrwkIpuuvRyYj
ueKP6C7FzPyKGL6e3ufw5TdhgSMco1R27D9cYnKobH9eBWY43CaThSxaI/NmbKy+M+9KcNxmYGrP
yV7ybhiJnFhUFhj5z9lVN3MOJfCASLP+j3r85aPHawYlO57RpY5rTZeKgmAUlYNGlvpslyW67aoU
Rbs0UM5wi3WztvjYLkkUC1+oTfy90YecP90qyGdFmIsTFFNr8F6ateXbNwALCuaXwo8+FXD+gLjT
/1O0oC7Q2F7xVA8dan+HTM2yWW2VV7QWUn2SIAT9i2Nua/Vj6yaS8JWJdnTh/MEfNUnS2QW8/sMp
cUiBaTaqtF12j1T9P2T1s2hfocq8bqqw4ZS5/AMwhMc0JMNclBDLw2npbioM24FSav697CNWpBCV
SBjdtOHt750JDfjvcxf62E5uPbAw5zdi1aN5OMmOE1k+3KBbuIZDYpzfXnYSORiufzvUzpmjNJ0+
W9TYL9LG9YpgCulh11AZequ5eYaHcAPBm72mnKdEMzsj2IH8JCiCy98/wAwLeCfVgyqu2af+pNJU
W9Xhu51PJyKGQYb3BxpP7F/gg7nDDVsCj5UypZhCD1mFStq6/4OM19DspbC+J1e5Y+Sos7NNzqYg
QwOPTDRRiVnDuyVz5qdS2j4HTtrknibI9SnMVIn0zM8fHps0q4pCqWVj270scRHYAeGBmcA3XhcE
F/q/Q6rmyuNPmXBIE1BZSCA7vx9YQMxTiLrZxxm8hvZm0nXL3l4FA9livLr+n5Cn5Nw2/Ex3rozF
eYRQGocGYW/bbzPkI4VLSWsVeIjOGGhDOdzjXqUofX4L8ALQJ9ECUcrFMCMYahU3oaF+025wLbAt
rM4yUdpK1kckcUHpfDpioISKwfNE+F7UpU6/UYFrPKUx4pn/GV0noN5XrNDU2c4lsV3p9wvy+ENo
QZsNpAau8+wjGJ7NAY/dKKHkf43MXo1JYb8hdI1HbMsC3DBIar01zH5dPVEXn0UAmznrlb30A95X
OxnBcY3aODcMAdD75T0W4r8ga+tT7axoishu8i2LhlCzs4IoZ3TpVx8jde0DLlFCY4tcJJFPMmhh
3s7B3ObkFMa2Mwv1y52Ni9cUCYExoTG3IW1WQSp5Nt0PUAHxfDilYKvIDa5WymhQVQRUEpRJzhIt
9LzG9ixvTQrciRwQY3fiH0l+HENzOYeHeudGt1DdMQkV1O2DE4T85NdC5Q9AK/OJBQy3m1PlHXG1
emIlTq0fi1nn5AbCQMMCD4PbGKwHIlIGZtjvdwG4F9VynbNmGwMzVz+kyOaPXzFtTeEj0yg4CcdF
z8DjuYgRoFxyamQKgsuPLkgkpx54R+UtnqK2wXA1Z3BS0h2sTaoKVOhgpUDIYzzcz7auMdQDnBwZ
RuL5lvNySlxexoehh6j7zCU+t2WiIpawNV1Rqf8rLlZqbq8Zt7szJ0nacQ0sPCVVAY4h/GXagbo9
SosYpSwuIY+/2HJnJFKA+FvXxjg/ZI1AEprSd9ZXIEauv+usr8r4w/X01i2fh275bveZ8A4SI7Au
REjdKegvS4mxVRcb5C9BDn7qpM3R7NUmrrti24xdYVnCtPFeRZUumugVwiTI3FvROnQ0mDoUUYVD
R8sv25uaMEeSrtvwu4taywTcJHxP2SKGsxFOVKOTL/tA7prso2eiYfGGb9WZM1X9hfNSrSNMhMnC
d5aOPMi3PJ3vfoPT7NgrrNKreAn10DgMWOS21NLbcJDKEuAhaNVlAZjpJc1hazyLoNmRs1xNTyHZ
B9vJPrUuwxc5IUU9LZbkE4Fnh9Z/UDw5CZx0yEW9iMAXdAUfEjBrUAnlfFI+MVwfG7ImAbip7dPe
AyfJf3gY7QZnd3MFqYDp6LQjeBDnJHlQ5JTwIS1+DatlEfwMMnYPH2genzxbYgsZCihivOT2pbUq
XdodsVDFofh9BloJDzPuq3vVRC0qdrmyGiAMjCVDQ+PXwI9HXTjAZhoyoabYmkI78fkNJLnWget7
BE9bW1GzXUSZdbCg17AGMFOZTgvdglLNweKm6qRDzQozttdXjrHRmiZEeyNjcnv3OwYnHdr/J/Ms
1arLVLUaXrJa77sfApZIA36GaZoNhb9M1i7G5hYwN++87Lrf7BNKB0y4DYEvM57xVNESMz0tVTNM
fpCJHj0wE0rvMLMtAbK4UskuziV3r7fGcJ0mzmIlun6GsEtkLKYhGZMf42DRFwdNsE6spJVXGrJf
VWTUqhGlbaKM1N3PBrNDv/BvCbL9thAgTvgwJ2Fs/r7dsp5q1o2IeMIWl32N9YdElFlQwVT9rTRT
A1TMM+ifN6E4HJjKcHf9l6svJyru9swTcblutWTyqIXOZTyT5pQh0fku299ZaNXI6vpUzJnJBsUd
OzoFYVgrug26ws7b3mJiZ63GiCCxjq7QV3AcRAEU8uqP9H7DO7aUs0BTXfFTGlfu8pCewZkU9LdH
5xH5b/F4V2zhJSNo24o5z2ElAjQK9FRWcNvqnfA/0p7ZW7LaD8Rb4O0U1oXVrJ6LkoLUx57u8Uzu
8W3FCgXLa7wSrwWo8PK9qeyJjnb4No2fhGmYaYDPpMKKaH7S2cv+LnmARRp+dXBQIiJXAAHG8ITq
/y+oVKb3ZvspVtmzGwXBH7gMVQX2rEDa/IieADeueMAutKX3gJKyVpUgap8p9B93SgeMcEKt0Be/
mKQOELW9Wzufd9RTGARmLLMBse/dDl3ONbQpTvcNtuP1ijMr8a/egCbSyMTheBKfv5GbBE6IpAIt
S40IwmhSLQ1gXpjTdDZzrt5+O5/6WLi/E7W+/R4GcxpIfd090fYN12s8Ycwf9t5vvuOpsPzF2/1m
wzPnhqw0LJeZHflCzaW9c13N4e067YF+0KGYHtMT1LcWlsliVX9V3DsgGnClkFcqG1hE9uqzk3AY
gn/5Ft57/cNVunB/mxO94SYkSwCHW7Ijpw02NgpUQmr4TV6MjxeW9bZiVrjXfwhU7ZJ1Q83i5dGf
f45IlN1rCjx2pjaedKKBTKbVek/o5rYZmFeeFx4K+yPLpclO1GwPZPwQJVlQApYZoydqaZIanLhj
+0VKkh2Cdhrbe+RHZNSnN/667CFekOdddXzjZeCndlcwIm33NUFBgI6g3Da3GcW8Nq4cTx3G64Gd
cEwr+Xvp/rHoNY2yZ1Eszad6FZGThJW6zySTb2oC+Xu8zkxKuh/QLeKmojvd+uAKffhwaB+xsKnj
VsqAvew/zz2oxxNrF+T+QN39Q46CMMvsFDIbOXvat/Hl0ELhFlWxHTs1QjfCZh2R+OrilVoGZU4j
KPBabekV00pPvESconZVL/6UyRCnsnHovrQdtgy3mIvjwWv8jz58TaOFgp3wFV5xzCf/+gcbD5vc
GeRs9gLlTO3Penonkvxh3b6cmcdxvowrRWVXq9w2pybe2dOHYtlRB8jH1Rsi/uKwHm6cunChtN/x
SpVYAJ6LuomJ8eFq1SXn3GLTPaPLjU/uRBDE/4pde6ImLioJ8x+7YRm/fW/ZeG8HceLIilJL6/Ig
O9v0PhTZtdkceQTQQfb5vh9WzpE6E8mcpqVv+9Di6QjmjnMzsH102ziDWm89VMV+kdRgazDIgqFw
4s/o6R0mfHoR40sshQbAJ73SkP0zNqEc3KGxgLJmLcvSfeci1GG/yosVJz7Bxmpqgt1RlLazbSFi
BLfkSyyHuOjQCDCHEMqeXq1w
`pragma protect end_protected
