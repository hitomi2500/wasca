// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Klaivz8UsqZ4GOu0+R2sk18CsSjC68fvlyYqIfPBvhr6F6kYR3MNrbGK5mnA+yScsqVYvZrws8QG
Chk0rpQjDCmwHrTYCY3olNZF6V+1118HQs2gKUSNsyhZOdsfsUMPDV7zEspzQD43d6V3nVLqBGk1
T0vVKYhCWU8FOgzLFCJ5dMHcCzZdWkiIalG3rMkofB3Myfn1AWvxEBR/C4vYd036IEs+4RZDCaAj
rfk2NQoIA6IhQ4zP2PG8sPqmtzAy7IYnp1rf7FKoHuRwrI8DNziCuboaBkJu6WIM11fkhQgFg0/I
TCnivf2hUkZh79fP7g1RwVr+s+CtVCNdeAJ4zA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8rUNxUrxiyWP858BseVqV7kwhjwhD6eQ5NGmFk//KOTyAR3HMCaCUJvpBXltPxm/ZwN7AK3v/H8w
TscHbkQJxCKxvcgIrDfunbtNZFdZMPdGArpWzNcvrtuj7g0Z3HkZGR2/p9Nxf3ioQQmQbDEfn+5s
AzuH9YywmX00J8uA7XNPjtjMCjI2LCXMafURlK+ZhthHB1TtRV/BZ68bMZ6oSK4z0SKX/n783tV2
TYyjsg4Inf/kLk65XZQ3Tz7kYunHp7DGCWS4UiMqe2DegVSkhvmysCZYIG9/wBRgk7nnC8HjQybE
Y8IBi7NrE7Ns3VA0ZDhXrjGtRTWunySEsERWyb8QCGPw+zbEQdwH5gag/eM9lVNU3ZLJzwq7/9RE
jplHM3uq8VVq+vRLEgMeqVfvj5bcI0R3H+Vv9szrgh1H8mye0Rl0CeCmVG3A/RSKGFyUKhdmLx9o
AJSh5M2Egh7Q8djXDOd4836MKcg8iGVuIvYju159dUC4NQh0lfTKfhal7G93GjLfTO27f4o6RoXR
EsfJ3ll9IulwkxU7lH6syBpFOUQzXZF2TfGjEVbRqrSML9HHyrS8dCyMzLUTaZzAYz/nbNrF3lUP
o9tJv3WS2vSzQPC+TCUEMePfNDLnxl97pGiZg3UiDu6r4FN11ON4YSCwOukqCGA0Xoe+vhW96TsZ
C4laCTZJrifR4TeCXxzNB0PPpTAQMKK/G2ZUPO7S81LihvF813Z4Hell3iVREARtMD2wgzmobtVc
aViMQFJhVlQYefUYgmTojAfXK5N0CB1Ue8KOgzp1ukL7jeASEuqGrJ4zUeRKaPl3OSvxn6OIMu+V
tTkVh2oBpVIGWtQUwt1tDyWeUivd4Wmuai9LPzY63oBSeTDPP8K4RskYvoW3/6WiCP1Y1HFmt/nS
Q/5YGgjJMMvxzAn1Fgt3pjFON8Pp13AzX/t8a/yW+avh2UN0hHz0Y8glGigiGZwP8oBXuvH/9xIq
vxzxZvWLDv4+7iku+rdAo5XJJ7NKJopK2F16NtOWhhLYqXGIKs5gzl2gvsTu255C5wuwuz1hfsis
z1RnWfgCDPeDVrWiEkcbn8IbWqsI3/VN6/+dRFiRq5vKwK5gmeeU6nS5o32r7w3kodUBrgVjWUZP
P9XNj/ysgLAL0UeE40frvkNdGVzp1RaPn/Btfa091xicTkKyHI4ws/gktJ4piCb2y2RL7PN7PQTg
qYzEqN99wpSWpLlhcod5GVnrWRqrdD0BkIxKkHbRXHQvhsAXlS/F8Yd8Fzo9T+pkBg3eRylmmHzH
cs6LfaoVByBLiYorC4IyZItrVV3wfd8KhItw261nffTEz/TgIPUsBzUj74EUQRW6yFnNBaAOOmR5
T1Gf05nwcZ4NwgCICJiFrUiwSXoN39JJ1GM4BXj5kHCwvBmNMzRDkACRH6E+XqAe6g4fX3t0r5y6
fhR+/cpu7kvN3SPjzyZnNfRn0UtzX/Gf02QF+zzlpXxZfZHa78m9kkMteR7O6U8A41pznAFyDMoc
OnDj3MsuYhZuegh///eA50RfkPs0Z0o6xsLAwDZ/3AfqrI0r3EqlcMla6TV9dbGmJACiN81uoGoB
Lzhmx2j2MF+uXcmBFm45e8RhN5bHyg1GT69Z8v6ttze4Mz5UEB8gH7pjyGjujG83/8y/qHUfX9YQ
5F6SpTX/jfX+GuCjnGXr7UjMDp2wQnizzBLaFINxhFyO9Ku9W/+Bn6ZLGG3qKLreYAFkxwlk7+cJ
dzIgq5bnCuJ/AO6OK0X6HZtuUPG8V+H+RwthMJXkf6RRQyYe81OJflIZtSnQqOygerhm012GTb6N
xZnDVSMbtyAzj08Tlv9gKSf0V+hH3CwiNdW/+nr3M0hgY2RQQABMZvsHUypX1JjXsDRasZ6Q1yU+
p7FyHiT7UTBuePiAxj7fbOVeRNN7hCoDyVq/+fba75PuV9gJb+cr5M0IIWYLCTK5Szcf4Qpm1sHy
UQ0da+7vPGpYQ46zut5IKaFzVluv1amvZVyoq/fMFgqN0TupJW4fcVrNppXrkF7J9YnPRVmbXcQf
rKz9BlidLze11F7BVJnAOBvAnHTV0lFIFzn5/UUZoRaARuGpdJMcb5qRV4qRo0pM8BK+UC3A5hAg
OCMZxGrXZkFMeJ0Zo6A46loxf85/IjnI59xtZ8AOupdyvp7wG+/e1oFS7ojRHG2Pp0PC1rh7kfS3
K2rMfCqW6Pjg5wtwLFn2BmzSrJXhwBTuoRv1int1ikoBTsDSSbknyHr0bqYviM9/yWTQcZmfACuw
Gv5g7l7L46sd2Oe6n2f2N7Qe0XALJ17nwgxNXTPNjYLP3UGOfqz0vHO6xCqfc4LhvVnQml5wxIBB
XKtKl4PpROI2ge18EOhcm60u5Gmh3rHYu19PSEcvsjso4aivuK9gsArJA6u05ywroZlKJlyPvIJ1
CATuvFpF6zTEgK5rXWbJLo/3zGSAh1QmisQdbQ0luTDJ+yYppCkGrzJJ466loxDc31vNBHy34QJX
QM1Rqp2uh118Qgru/BvhYNsqw/tj2d1nS7vMTAUzpX1K5SxR2vjVJvhLHGyMCEa9nZ0wgjnfY42/
+bhuX2fmfqI8T5roQNOi1wch1GZntaT+fRDjAFm4+vKVEJSjfl/j54LdfJSir41ABb6mdCVdQ2qh
/p5sSf+G9aieB9S+VoM6/6k05dizA8lTEbHhJbUrNdoiqKJfcM481Xah7h4stWMc3p9o6TglvstO
n09iE9Zq322zz8aXXrmNMkzgC+/cStaDOxTQYfMA/Ack8NDYntTaK/st13CyK29JwPcAjx2RfZ4e
fqLHzxRwFhkjAJnXSW03VoL8hRlrdTLmd2Jlrbt9FcMhhJXNTe9ZDwIO1S2nz6vAgbLk10652/a2
Cv9qccyzAYfFewiiDNXaSu6f99lCeCHya+RQ2JWPkHcII3tmbxceMxdLy0KYuvvRFApjvoWK6OLC
+6rsetcBsqs3SONaajPqnPfMGRgOO8na9PrWmvCC9GXSYYq6GU4rWX1oi9Ym+mnCheUH6tBPDmEx
35ch4OMCDJQZQuNCATgcruyFrMJ4RuG6sxS4TkXgBuL5k4SyiddsKzvikT4E39b+57LE92XSkX1u
3TeGktzZcJIZvWIOlaQbAgmKPOcKDy9NnigAiM1gmRADLuLbTJza1HFIKPn435XvSEmFkPGArOfW
EV8An1GO8q7r35+RbhFw9Ybjd5GDFQoNtcxb/nzjqd7eOupz9mSfDEQ/gMo0dkcUp83ZpeiFDBFX
uIHyi6tOotH644xnNJdC2LTpEJ6AD9/cKV7Vyb40xR51n4pY3+xBqljmu1i9J54DqzuJSlzuPk+c
jc93b+I2kCXkZrfAX9SHq0FOiNuSD/ensAflfLT7clPbtEflVhj3bKCIjhbdrEWCY2Bwf+J1fls5
5XBY680XgfhGok0egcJjEINxkMx0EhZ+ktH8OuQm0PZWV97Z3mEnZmQTYufohEKpVF7iZJaGI24i
JygJie70BhKnYvQnvHjOgNKaRdSXDhrQILHntBxB97PxjT4GFo67B7B1Lm+RQWnZ+CNT5iWuGHTJ
/+5qTbTdCcTmoglF+66bjvMRIXhkg72zwIvDUf8t9B/4A4Xbctazktx9AZOXoFBtQ5hqWB9RdkKc
AymnIHkQdHlAvW66iMLhooa9M0UUXHDQkHl9vS1a42vRPCdbfNELpHw3ONr5A5uXItWqU+9Er7zy
rD5llw/MwInTqO+RJXoAPQYNxumyO7PskJXm7is6vCQpI2PKRE5TpjbfL7gmRCEAnAI4kKm1AA5G
1yH8kCLHc/18Q4OsoGpgzdv0Y7DvMEcSAEDBKMOOXmXq/4K7KFtXQGRFNaW02YyakFLkK4Gyf4F6
k3MFcEUwt0qvI+8D42qmTHlaTTWrhBor8nm8FwtN/8iYdUKsiRaEfvtonC6kpx7kqt22dSgqhz1D
4vNdkWlQD7Tm8Ul7McQ9spkBlb/jNCPq4ESQKXfOcA4OcaoY2rjFNcXOklLEX1kMigqKKZ0kWQfZ
ERLjSSBZZOENSoBR37j4JOIpys42kuhmOx5slaZOqGNl+siCxys3IqetKhstDqcMobJxGkhJHvQ1
uU8HDW9Ww7RlXBecPxsa5PAhGnrZBwDn3rhEyrsXmohe9RA6e7rUrSfKCNwBbdMQxWJe00Nmmhu5
8d618fXrYyEfCa62jT4LN5ZFPyTdcq6Q6svDBhne5LUk6KxbiTCrJ5bBWxKJx1mIBt0DZH3Ru7el
CopbZ2Qb3ZReDriD/yXgbc5wdimqaVhoV8KsPjLhRvGWCv1DNL31fwKA7Xrqul7MGDsrTza71yfz
MgNjBh1PLlVPxuRovfKqMPrW7u84tl0/S6snQkgt+xqQJSCxQNvRnVLqazakrG2Ap7sY/6hJAgTp
xN0OlTfnSJ+ntYhNSW6x+Ve6oJSlUWtm06gp6LZeuj+BQbAOZ1c8ySQ+YAJ7bykrs1AmLKTdJqU7
9qZrbfV7uxr2k9omvmi5C7faW3eUjE68vVXdhSuCT1+aiPqRN0kOs0ETaSc/W2uovlW+Xax83YKg
CdPHpxpM+kTzKODSlIhHRJXxTHGu86d9qj5k09V1+mtt657atpZgILuZ+o9J0PtzP2TYeb6fVTE7
QN8AwOOCSsLeAD5XU4jPKlrTYleucdD1ai/F/XRJu7Df4AuBiPgNeyPbttAXlvo3YIEh8I6HdwsY
8+FDqbaHYhe38ajB/aehQP3Tyd8dGHM3B4iW7aeLQwaNue1ulHXTfhoasqatde0hGLFSncCS5wwS
J6YJtnTriAS1Bbc3MCqHCi6RgsEC9xvx6weRZ/0uesE3mayBoIBR7VSUJ42hiBGx1e1vf0x5t3k6
o+Ar3kdAwEmwzEFH9GT6x0TlLHu9055iyv0f+4OzoUXC21C3bku/4TKAC5b0iWoLjqUPFdcX4LES
8T/Nm1SU1xRl9QVPv5fxWdRFuyjWVW2KYNcmkAsVfcuRSBfc1br1/f8wyXUOAF3c3P7FZLQpE5Er
0M+yf0yfJCdvMSCW3zTG2QF0wNlx0jBKvVDttP/Er6H2DoeibHwp1Edq4Zq1l2icZHqYh85gplVe
TbJpvopC74fM1FhyDYibxyunqn8F+HQnxUhdAI80b91OsYHh3CQ9H3b8XmHgdTE+pXehW53m37KQ
JLYI4woblnzjBeShQ0+sF6UmlzfJ4jwFAL+Tmz2z67VYbP6X23eZduCBV3kd9si7GDD+uq1V66z/
WQGZ/kwmQ/0zqM2bvvLfBM8tQvbFtb8SMNyBWpPcbhVxZTc9KD1vCfjkCLnriZtTOEMNAQoaOG++
FXwyY++qVQ0bEx+UP2Czjpf7qvM6JoEtfSPgEIbbaroBSpC3KVLQvET5TIqxbuBmM1u9PFRdUtF3
Au+aekttjqUfr244cunc7dd/kfRgoINS+CSb1eharN1GKgIm7NEXiQe9sdIJFQ8DpchV2DAOBWCH
d1oQNYkSGUamQVXUvpCZr2hVzN29b/++JtXP6tI/cm6sOX7uA4hcXJNdxwbdk4ZlSnBXFIQntJ1D
q7hX0rDQ8Wjc13WxpP+iuudm5QFQwb07lJU5igts83uYM8tNqqN4oKIV/KSluz7guL4VkFTyz5ZP
cE56elUTGUD/If4lfpnj9XY3+3Oo3ENveNEJPusoOSMuvNzMaLvBaZ1+By4fUg6s3NUfSeCWEMmH
GJxJzb8trHq5jbszmxnQ3bqHLi7k3QS6e03TNz0VAqKOwcFtrHulYSeiJnxQ+yfbe+mZQnwGzhzJ
B5GKzrlCsqZIK8Miub1GGrBS6EdLj+MUkAg0lLu4VKtyNJ9aP71crbPd5btns0CD4anVIKrX3iin
PFFdXMZTIdBwyXxiH95LaJsI66OBS1ErR6wJ4/BLbYnksGDmmCJcp9d+tZaXa7/Q+5ahYEpMmQSc
xZohFiR/R7rjD4SSNjeQ23eg7TUoxUdOSLSjeetN+rcb1MjgWYD/DxzXWTCwq16QqfdrtwAe1NWF
5ClZLNPdVmUAo/4YtXafVQL+kOktzK+xUHJaIqsA4Fm2FEnz4topag23tNYzgLdMGBHVnP7Oi0ck
JNcYbxad29gqEoQwH8ANY2NCHdC917oRBOZ92jC9pYgR8eu2871WTH7n6hez73bGfrcaGViTZZHn
d0mqnyJ1guWMXw8FfIZZPirIEHFAjux3iJdy/YpuYjcVItG0TsGIgDkp7hJ4Hp9ylOcTm5QrHDaX
M5+t5cxuHfBzHtR3Fe7vd+JEqPtjucpxaHHCl3rqjghpjF5CK0Ew//Mwh77oNRb1PNUk+IDqJL2g
RtUu6VZpZJgVe39yvBHErM2Z8UJfClY75h3acHSVjNWeE6MEOShE9cOjZmcFne7ZdrjpSwimDUxJ
BKIWD5JiR/IUnTNKL5alUy666ZAh7sVK/yNmXJzksANFpIm+nn6Ad1KZ1NLjgh/rYvq0uonWHueI
AtePqnt71eAZ31dw1A3ljzVx/sldltgDXd2I3GtsckaNjN4cL+FoWaP5oj6XDnZZhQRqsC2LLKTv
dg8BjnXwMk6F8vVxGoD/sbKlcDRWTD6e/huf0x7uqr7phaGSxWUF3cZFM55ZEYWm0oarIf85oALi
bK5f/ddB6A0u1PH4vbex+hlmdq9zN/gXuHR2Dxp5s6KpH7BKg9k7xN9P10ifqct3uMRbILZHl3Y+
XFgH+3Sy91odx8MKR8/INnoyPqgIOdGvG/ObUvq+7jFl9kCkCm0qa8lJax5N2Hkmd5HcBKVp8EmF
lFsYf2dCEcQzMgTPwVUGDBNbFXdsMdWE3mPZWkQKzkVkxDDFTGOjHbKwYhmXIatzC6XG6cG+BzOB
0MTrDaJ7m/JI0HDLaeM/M+ir+xKEPstkK/7zIWGDOzdd9yKW4uc3X8J2OnhMASVvuAGtLe3AU8DS
n0S2ms0cDK3RhU2kfPVns1UNf3OfVIglMNUT2Bs5SUOBaOlGOYCccSvVXU3KEo/w6D2dG8s4zF9p
MmU/qwaoOe2/vRkiiV+9s+Gobxj5jb49gE3UF8RI07OIsFxi8i4e30BMQ6Ex8IaSsCGjAezsdkmF
fhZaATkH9ZLWfCreb/mx/J8ymPk2qkXFpMDQygPcHBMeiyKVI3xexKc0bEs9Hm68avi2mrLv7M0h
4NlqjQL8O5j5tq5VKD0NOKUQh/FnFgk24M5zNp0q2vZ6CxqxdEQruGIHD0Ihr8dekgFIBWJR/X54
GD4C2SYXCcP8jha8GqpZ1iqDga9KoOXonFej2QCkOwTvGQ53+zEcaVpF+tZEL+AmjfdmalEYFWTa
yf38Ge8/zhwtznQ7G2dJczlqqUem2I6fk73ObGnl287PnTc9HbXxVvikdZK4jd/q50twHKw3DzRg
qIttNQdqbVNdEEtHpaXHpsKfl2b6B73fYw3eVjGK+ejL9Lo0B/tO4KCe7SYKgw0vh55DJaDtuvyN
VBy8O+XmKCwfpCqAg9F/K6Y650UJCg31cPSQfNwGRwTvl/kJhbTRaQ345DV4SL8QcthAY5AcZPIJ
Y42mUDiB8Ue9LD+ww0nNJpWBWHZKZWvxkhtTBRoFuM8kZPASKCRpmvDpgYKaf1XFQD2mXkIqzcXy
CPttjvmSGKecW6+JR9qlceXSn3hfc9kNXbEjp5S1JRUyRSZ6d4E9nISiIBwpCvB1gQg+chxY0hTY
S8rT1CvWrxwPoy2+1yuzcYiS5Y0hiKVFl+KIGt3bdn98OvP8eEuoohi54ZuyWsc1TvL0c02fcmvv
PEBpKOQpGZvP7ECLcalYC8c/+yHYnzD7ddGPE+jc3GicfRBkyMNcW6v4kWGCfR+SMs744rJN4qrQ
2sd9UQB6wYR5WSI113w63vA0qmi2YTzYbmJPQKOGZvRuopDmz2wNzC/0Z3SdOi+NQqsD13O65GsH
rXHVA5+gLWm34tb2CUxizQRNqRD0APKfHy560LMyWU3D5ISrnt7mtSES2M/hJORWJUP6jcRaztPA
DcidXnY6c11xNo9gMsEceLkbXX4jP/F9enYIk1d9MqVXYa3X99e8nsgUpEmWbYDJKH55hlD40Ytj
IZ9EAgJSK9paWiYXJbijXWxvtrDVd9OFd57RkTjvX52seSAv5q5G+N13ix2QAhTmEWGxkAcVNuEh
A82ReciV69zdaiAKyQhZG+VAqQbx8fx7NKOELJvpaliYTXArzU+ncymkY9+pveYdDQosJjbjKsnB
ndaJR4WYseyhU8dTs6dg493Ao5GAKb7MMjsCJhv92hcJQDXvGoSU4VChbBjAYRTUgXS25mc8EGj2
F2CtaGfL5dArAKyoV50Zx2VDXRSLAxq0q8tCjzaPQ1jJAwGS7B6eeJ4P9Nxa0rvbYspRH8kTXsoA
8hPSB2LIQgcNBrOO4XKkQ/kkOhMyG4NG35WZt6JEF2IdBWUGG65KVOYnd1NLpdSjd/iYtjymtg/v
Ws3Hcrw3A9CSIp7YGfA3MYVdzLpnMMYb7nBTBdwjnXieidkRYxrvMT4ZC6xyfVycq+Q3pLQ+RiHa
UZQuKWXmIXH9af4ouquvtjbRrTB9h3YgUx+HfI9Q+GGvvWIwzCDjSxHe6qUT0aD0MNsEpkGGfGNy
/4gICsmyUoJGlGX/MY9KB/NcwK35zKBNsv+mMEfcSc8mlDDdEXXHA2rQQ+uIga9LClWQNI/fPo6I
kDGTAnJWTs9sy/bqr9SeYBItT/bc1qlC5cBZYqq3u25XDz5i9Y26MM7YSIF/LGGVkioDqrNpxxS5
+egyFKdtjqMp7VtC76y4avkzvZt0F5Rn7FVmS0afmc4M4MnkzRUWzB44Kx+K3mCNpxkzTSfc5Fhj
NBdyV80qc5kpWoIKyNVTV7zi44XtxJr1aV0V9XJeN1FrfMFJBQHifq9N/AvFFq4DpfntN/BaKAHC
47svv5nc9Tp8nAgvZV4eqkl/0HzOHMqYTsNkz938OJTiM5jfxAEVR/cwWijg9drYyvNd72XnI1dn
CGd2xcKRDsr0mXxSY1b8tlYyTdXQbSi4pvFXxIRYmw7YbgDXLt1fJIgOhFZjbZNLkQLcxT3X7+fc
GuW/0l8mKd/DESvfjXJoboFs4yaYPQQpAr5LaENjEQU85lDKmYBy2sbA86mARYjlBDsaEYAQqU9p
JsJjuOb/pxnPoeTmVQZft21FSYD4yjHFId5JNwimIS3z13ooThjpk9cl8cm5vvW+PKc/meuc56Lv
iD1KKT4eivgAIhctVw8cN476v2V8Ojp2I2CKJrgN4JxCZkgDQNvMpsWCBndY4xNUsn32aiZxacmy
FYgVfAVErQdts6Q9FNsX2bNB/5vcCjwaOqneF9uoWXKwiufHlkQuvbIks0aOqAPk8lrwEMe4/oxw
18EvznRjVCVFvCcR2KgMVM3EcAb3TUzDuO2nU8sceXL37phu+PGFRhEdlyO33mdjsMAvEcLpeM1J
2fFm2gjxu9bf3SlbwogEsFvhNxF9h82/GCRmVQtfPlaovPL0kO9BEypfdBhzu9LabrOuErMLVPBe
T8wHset7X70FuKJJj7woSQtKY+pJlRiDui0eMGIHCrI830U5FMmh/ZEkCwcA05rqIwk6HOQJ6aX9
hyRsZdWVlS5EtcXJMObZBY22dd4fBGpz/+PGSkKa9mzpNsEiLQwO3ZDb6q5syp5UImOkNZ6Sj4t1
hzcQuUBhySn2QBuw+LgwzkPyo86T36eSb9zLCYI6mjrEVgIJfJztBZLjaKCEV/XKXUqLy3oZM8La
ywUgL+818I2zt/j/yZBjULG3uyc4S8YptPkbW3H3hb/DF9p0uvCZXoD4FT3lkVKtqmpBkVxH/OJK
0raYCxZ6uDgCnLVoPygVLaobvnuhgTy/a7UApqbb0FkQANMEPtMdXnYHZgrVP5at4g5wx4FLlmkL
itPJeDu/wMPethp/nLqArs6ml8tn4E2bdJZaQ5NY6Xl8Mcu2QbIiTsI2lSqA1CM1c1N7PXFst7fg
ZMHE7ObDKEF9jyesncV4Bksf1h86bcfFaJ55Hjzf4SKh8j/5UHDFYSVfjtxWkUrocOJP1iD1AJG2
t0euKxpyYzFmEnpEBL5reP9IkIJMI3FuIsYo1ZHBZKF8JD0qbAj++CO4doMRoEmMMsZgu4Y8Ce2C
OVRzSLWo4oouYx2nRxUtjiCLPHMD1x5tj/5kLzfZOY9p61lqh3r+8/UZ5X7h0zpepkBX85lnES5k
MKGtxOd8MOsXzIgwmVcDINMLbBJWpPYz5H3e/ZdWOhsoaAl7l463/S3FMRECzBC1FJgqxz2sBOSx
R3rFw03+rZ7p2LcsEMl1oOjoxPo+cRYXBzqFSdB8pQrQmZWsrmRaqq1kUKOFADtBh0jeQOkDlkE6
Rkd8wMiAKRwF946d3+lSqi2WSILbJYD6DFRL9ewCQeMueiwsAZDPhCv5lbwWNUmIWz/KAhCsG7F8
UDB5Snced/hkBi8HlXW8Q68rxmMTuxEAnTLgL3LEXy0BrpOdkT599VeTpeEu2J8hjwnSXgtwQMQa
k7j4BhIn+ia9LuTky+gWvwWKU24b8TovHPqqiXgvsjCvhjW53RvWOHT1Bxt4TgoPSihG4j/Ye3QP
57nk2BMMdx0RbM0GGImGAXy/XVoUV7JgzHxDX1qfGcp4VoSwD0IpnMBypJmK4qGyKl01+U4Fg+lL
MmKY410N2t0QuTBxN0Wxu9CnyZvLE+wlIcrShBTo28EalJ1YRoHVHZjl480DABsajjkIQyYzjOHR
BRnEk14BjF2edfzf6LkK3fVh1syfkGT7dr8QDfxZiXnW1kN7jpPVBSaIiuugVP+rBB/d0mSvM72f
B1hWqDTVS6FmQT7JsR9L9Na4oKw7RojfSfNSFkR8He7anQ4Z5ZhH6s5xx5fWNYBf8ITFVJqNVC1X
02xRu80gTfwtUv0qQKoebZEm4TFtJlT5X1wWX1HRerfoipiAlqij4O9KoWyYvgfJjoZNa0wnXSgJ
RoHPMi8+p6sEpRfzmwyqEccpcpjhtWLZd+er8goaRnHmit3jd/zBCPNhQDQXJCe/y7ck1feowyPV
HzyR/YpU75yNqUjFW0iVYrts18hHwUQsrO0GtgdZ9coqja0iugWZEBHQAmBEgL7/EQbHa5O1V4tk
XDxXKMLdx6nun6X3ltP3CcBsNbjsqRlXe8npCMqfeKzfIShUaiVE81IpwxDo4T+g1b5NamLmBtTx
jltJ6dhsUvXI84yQuw4bskymJF+Kdt82HXj+Rj2H4l4nuEYbOBV2Ax/NiUTCVctHnGa/h6mozZJe
f0el209Trbi+z4++mFsAzF+9mjKPuwQN2/MWcBIO+rW1EU1rl1EoQ8fs91aUsoK3P6WnV8Hl8mvF
NgzF+q1W6kdKU548Kdyzni2+RlqY6cYS8CD+Citng2IlXAF7+n9XtgP7S0SsrYbiQmbmuvWScq/k
ABBKLN1Mr7ueUjXtMRCyq1efYJWoaGTVlgV+BHwWF5tI1GFriwx4FgQCeswO5yw1aj8v1ITItzWk
XEXRiBbmVCQui8F/t/GrHmEc3/xZAQ2iUuIjluvjWJYcB6Y2EvFUCXs+KrU6UmZGHNdciheEXqlw
ruSdjXsHwbC3bdSkhyXpDvAWw+eJx/kmCFGdp0MAB12o89aYu7fa36So4eTsZjn8HdC0OBLbdfm2
xRsO3CvL7Gdq4YdQZHHUk3W5ftGLpmuMglFB9ExBYcw6M93ZL21m0Jk+wKWWnlGlunjAnKnOBHas
6bKtWtiDUx3LQ3mD7gjRLBrPfVA9mWHQsITi/qNCHFMSrcQVb4jFykfpDEydztFJ8ab99rTe8vSp
STrYVnOEelskuWNE/e5skTSY15OwsekNedPzq2X2DHprdYLkGXATeNERPOwH7v05/ZaWbYn2tJmi
vLm3OkAzXnz4NzrykfnwJ6nn7URoNQCsLM/hZFmHtEI9ofOCsSEX1guW7K+eu9rUa0GBzb4C310P
YcMl0T6IQdzJHEssPSSWekvY5Vm3TZeoW1++RcGAuXmhkalMFD490gxB8/ZZ/hehiiMw0piu8d2b
wtgNZbm2oF7OhrdvbW9V6DeRtJryUN63kY7EikcaUt4N/Iru3RQinrSkVj/SP3Ph664VMHqRLOug
yTJJ+0HkNvnY1aqsYm8o8xb/OVfNZpNhWOoMxHUFQmt+bhyoF0TXDR4AwQDERfdJEaZe3ZznJTCx
2dHvGPP+QEAG2foVUjQ8UNXMpB3DK74F1TP7QIASwX8miqatqSbWOCh++zPbgkWRRtVtY3soPZnt
TJQjrxaEhnYf40P6czSnTVt2ZETBmFVEcYV3OMMRQRE0J0RKBpz6g5d1fbh6+YZOcVDHBCb09Rfh
2YL9buc0zQhRzNc10oe5OEaCPdqJiZDN//oF9U5PykYJq7tUAg0PiN3hmXntJN1ks5Ozj/RZBavD
4bRtzKy+ZZOosBYbj/1CRR9EkUUu8LJr3HXA6FMjdDUnK7bvxVlI1sxK+9LbERvYe00sGt6kLLxB
M9G+n6H5Loq/WMzKVNz4SlrFeH8GEfMSy0QHLpy0SgDaEzPCQNApLY8WxUF7DgTAg/xDlm3a1aid
JwA8B8gK380Er04fgulL8xFNRpwsEkLafa3O5/9LLjfEW5rAlorhYWpht/p4DoRAF7cZC59bqaGG
DD1HWMHiGZ8r1Pec/NCPmDprBnI5LtmnmTEeN5hc1e3lVfer32fFTYSagR4frkNsBxTwRvrpwUr1
T/NQ9I35AMUBjkZIoHGfOw+gvNnwPLZUGXKg6pCcG9HYdVzSXyq4kgbfjpfwDEyBWmqJ83s/QzI8
hWXSn/Wk3Ftt7MrUNZIQfhjhL/QUe/FGTEIzV4Lqj1UNABNYZ951pQw50zKOwo+j7YbgwpLWuQAs
zCbRpLdU0bbYYzwmuSRImeLDnDn4Kt729rlr0IB6+9UCZW53nmiZzWmPgjSi7hfOaAl8jXryO1Xl
49CdSzPWRhbHNrsudtcZ0E2+KJDA/CC6c3pz4LInFFHXpC7ZxdCYNxxEcBXrG3gjUOsImSa5phKo
oka+4tO/uw2yFl2spDj0IZykugbLpGD+Z+m2P0PmxF72KGE25LAnBcYMwpqFZd7pR6Mdlmr6HjKs
bioVICz3yu5UGgUtIccGcPCU7Uh8LurTnmG+lHnNI22Zj7ZPyyL31VEgFviJRp/gcVVtUoD3DgKQ
R01xhwULrCgPX5qHraxU8zEM4ovxKdZyvXktbZ+v0j6Ub4DqGJ1OVikje7mJma/iESkcCkmyYqK7
sI4QFelaSabWH4eeb+oGLcAjxKjwphllcec/KPDh/qWSgvjhMdHgwrMIKZVUqevXN91XecuCGl2J
iEVzEFuckt5p73aaoTJK25aOgfxR8DjD/RzjJzzoR7HBRjsVByMJvBHOr4tyYgJNV9xTWeO9luMi
IfX7upp1A9u7mUhqAsIi8xhGeBA8SYoeyJARY8Pcjy+bfxnlBARVzbp/asBNNbMlh++1bXBY1tGp
eI0KwjkUlloMU/4F8J2rQOMT95iUO7ogi9xGjSw2+fAQlePMfYSLj/xyTcUrns2sCfczolMfWIX2
LiSzhvZ13LYKB6c8POHnlaga6s78Zu2ySmhg16MF7ywNDDntqKH8llhPnJK6jiH78JjAyQlGZUaV
nhBjfOYZeCy0wkHzN2tBETwlmDtkTD2JwhMLYPV6HW3src1eHse7htPN4kP0UjNU1Od5hIoJUQRM
/QqicmKwLLmbUiONssD5FdusTvpSZmWTGvYE3U8dWGqKAl2KlvOzjdFscOB8mfi3IBB2inUheozc
RrtPuiujzNDNoiP1Xy6jzDBRX4KFH6EF7J+diC0c/weOCMLzdotaEkE3mtCNwrXx1l/1XfSJeeWd
ovOGx+48klunLaacFO9SSwEBI3V3QwWO7DzkGbQ40HCFuUVo7w00J3Di3YWk6iNPniNLXsrnVcZy
Rmj6V5mRiY+gWh3gbsN7fTc3PtwKMxgr3QH1a0dgGxH4hhyh5ufLRTsGb4dve02gPIjoZRsPEEc1
kxWrmZRVYf+E5LLezxOg0YSAsPjaJoccpVNXErHkJBG5G9HTpq5IXPO6CgMIqal7vHD0Jm4eXE1d
uxelxCbtMe0e04orCMnKzAwElE/+O55O8+iqErInoSjHzVCDmjL9Zwh1H3X321FvFXJxZyGMrnUg
4Q0MUzINeuqUURnSGE7oQDbxVw95xS5QpW6wEapFjnWuK8gaq1OhVvgIW7N91DTs93iUh5me2NJJ
TlOrY4h3vQRPwkxnhmODB1byMpyrjqL3LB9Ayk5bxVkvXPi/Ed3dGnbrtpBQi6zzFBLA34r6qGed
su1rD0KvyCCl1V3fLJAa2yidMdzieytCyUQlaK3xUMsHMmprKWV0YF/yqmn5UtXICBy7/xnz5l8F
JtTZZ26CF3vUTHXQYZ2YZict9KSBmMjungGGYoOwfQ1ks8wcEqxndwZMH2ek2k+xWz/gxUOEFKl+
ZMy62OlAhdJyCVttl8CbUYOvoQUZGdgTDSqdjG06TWx4KEknJbJyCJmABQsY5LW0DKANt24O28UU
/5Uq9XstPs6maZWuqiFAQ/cCYv210pfg96t+17oNTQtJwkp6Jf61r11p/BZON0mx8RwXJfOeYeQt
kNfZQfgs4uXEd1aUoxeuSbHCr3jF1sohFRalBLNqkMjSRfHnQIzmUeF0VA6x8jqT8fEizC+b2GWC
dcGhrZHUT+LEjwLn9myZseUcYjg//5XnHKXQCEXAsCtKLKg6H9dS5T/IXjdxocC4J0ZYvMLmw8iV
V0wmIznRrTJs4ecsCY2fIKs6r6um02mgfxGoMMy87Qlnj+GH7gJcazLHOquYVo74AevvAC6elIV+
KlHVPsX8/A2eiJGCeqtlrXtNT29DgdTvJ/nSGbRgasbQeM08zZg7K1YIjCqeYHmwQrB1ZAR2SUHz
P2NhErJxF7vYnk8ZngleIKnq5bCB3DGArqLaZPYCWFRohhRWM0F6ztbD2fr1w/3Gj6PbYpGsXj74
MG3hRz6ZuCAdVNu1aKMItRlidwfLN5cMm6pqPOLtcRgSwOxCju+szHnF667ia9v6pStoENwZ/R6V
It7HkirYPtgBUNeOXwure8GXnO/qtmKTc6sDkPNYf5/ZHnSBRJGLcgKyKvoRT5dH7yopuzqWwRx8
hXNfyqOb8DNZXzEHQiviTeKf/f8F3yflDzquT+VnjsXeBrBLAuwpP7yx516pATvtq1qtpCzDTwCl
EaWFI55rwosjQHR2y9mBLuSEID5BvV4eTqLjRvPRP5fQGpucA3EJjSK5KXzY6BNNQRmzFG2cSYUm
8Bkwg8jkXDB5/c+ymKmXR2/O2GKgFHvL+MYQWIhabCS7Qa12U2bvq3ZRx3PPCJ8q1/71KLz1C0E5
iyTfO2wv9bPLHcxeSc3midbOZp2+06NUPApMvzFdlWCcWpcj1auJIKlxpVp+W4uUKKuOhg043KjP
9Ny2+66tpT+JfL6avv8OqULL4fTAN7W5VTwq+dl+XNH5vR5MK+CEccr7MKVHrTZ8qX4dFtBvi89q
F00jlRAEChjvmFVmKpzc1/01Sp88mIKgFNZv0kQGPKhCo/bzx1oLJdBThlCGRO76vDxEQ1QOHIa0
M8GYQzdKGDEdHcIjcG+5TNiptTnhZ43lRRPffakKgtxHjySMCHNLGW4c8yQnpie+M0FWu1Wz+KsL
/zSd8J0iC25frWPN65aQzF3s05/cYg6Kt86/X2MtCgAchC60AD9N2w8kntoh8Nr7LZCbDHC1ppeZ
ohFZLSfxnQTR1TWYTlfFGjWpL4l/H1E6I7okvXQAlmWekVy7RiAtKoBtKmtP2Pu5zvyvf03TC+vd
9ouvGtdFBxSqNT3UOg//eKBeT6q5DTRx3s/SINPoZYBhjRMIBsmCpQr2DX6rjsYILS0yxdTlsOWI
yo+/1Vqb2vSDpXDHYIvsaKiCiM+F2mtSwVwhHV6CQelCbldFI1UfieQFmOKnHBo3qCiChKdZDTnG
ghdmaDlkB9EOWvoMyKr6T4MbaZSUs8qXMCr/WSY95uRac/DcC30LbbfaaK/m/GdFb2p+O9rm8pI+
Rkb87+tUbQFJch++B73bK0WkclvEIvduh2iqtggFCX6QnkemHLyLhYxbi1r+czFp/j2ZIFyCeH6Y
fnGWoiMtqGdAS3D/Qjc6U95vR6FktNiFxKjZ6uzmd6nVAL+5vqLeha0PFn/b+g4+fp7cHYdI2+DI
MGN8Omml3inLEBXAD/aFz0NAs1knqXYy25mn8NbsLuvIR35RLWeVm+jQiNZdk5oF+FAUhdeVm1h+
uKIaESC/pYwjzh9N/dfC59t+KhNtwb+uS7njAA2CyVu7Gmmprd8pdJfSowUx7Z/ZLSJw0gmUPi5I
ZX/gJMaMmJU1Dtk+z0MQLLijvsQOyKx2AJvRQlkeiXg6kw0j4W747zh8gLpDrarar7O8gSNQTSsh
TABrqxVckVvNjZ8meO/YzJmG3pT15AhYDx/KxyghEq9I+TVbCCpBVoj7K45Ii8GwT0vPHDNYBjUj
4U4fhjWKfNxRcvKFZ3eXhNX79zI/xzuOzXYahHNTYFaQKd+36pnOiduuM/pNljEvVlnD4603+GjM
cEu33MwUGY28g1fF/sXk3ll4SovVmFWJXG8LmpouM4FLd3od3uc2IyT2DcRliKJGmNaymMNw+eK2
3zS4PM7XMgl5jsoiFHI+SAiIoChCWgRo3mtyAo04A15BCmJYYukER3c0WgSe9f4wZ3YApmHlZoez
I35M0j9bJbIloq8XtWPTU/5z6knpVycUuNEteGkgp3PLziecg6G9a8iyWFmZVxrXUWXJu2FVYLfN
GytHgR8Y+sOOzYGvzEqluOL6SPRyubMOaRSj4Md8l5etM82H+snsjysCzXel3f05mT8rs+0MrisO
iLlTpMq4H2cBwzTD+58Fkse71VVpYE5mpIKHLwng3bMf1KW24MsZXcY2zQSNhNjK8CSAXsiI8PZu
MSBTJM5pka/uOwJG41aYbqdwW6g3DWyzOze1p/gempauziudXslGm3zISye99eIPlPJX+Uvc7yeM
DfrPj1l18hYPcMeNVk6vpIz0M2lxP3M1U3+JgFPNvY1ylO4bg7Ouubi5hFf85CfwzJb7Cneiku/x
J/N9vBZfmcD8TgofpogDHE4vBd339+ff0UUDz8SBI6K2MjAlNYg8dcxTe0D6YlFej2JKi4bf3lSu
XAM8sMA+t38MnlQ6vlKidYJEReHbgy74+S4I0Nn0aq/+zn6LkaVcwsyH+DXLBwLBFEzm+urOmPn2
QV+pEgC2ApCi02COBouuogqhRK3IrP14M2Phqinh+wVYm8v5E8rFEHhPZppX2aRbGMu6brp8pvRe
tZn2eBnYhT0dUWTwC/BHjGzYoh5MSSYxnH3xvYg+jkI1qJtdYCdHCqXDXU52vVk9kHIo9W4FGvLa
rxtRaQtmKSwCKj6medf6yyJMMEw3EgZJyeLUJw213TBvj1hg/Ja1qfabKBuRMuU0Cf0nTO+F0IhU
Z9+jyjyBSBu4v68M11Mq0EgZS/pTH51hc/R9QhSIB26PlyU3a0wVyjoPcE2c4LXEAKI5ys2Zx+Mq
D+ePg3zmNfSZ2Bqnbv/c1TfKc7HdU0j9FD9sLADOLeSolipq6WJty2D8qGbfnPycFbq4ukWt15xP
KK5xX4pQr+ihRZM1DCwa/v+PhxgysakZUcjMs2ugtBcAmqNql/rQI+7lsiwyPquO3k8J6qzFDHZQ
4B2KChkWW4s7DXSGLpbczBfz3NCRbdclKKwi1KGDML+fAaV24I5YYHYUhHV09BV4xq7OAxSAnErv
KhEHqpIDQcG/jZAl1QtYtsH22CunuWEWbLrsBA/+t9HPBW19536hH9h6CU3BjwP7BtC6gJ5cN7ft
Z8lVNuwmHxy1x8MRXel1CwWlJm1ndyvfBfF1EmO3BudFy3TB/z0+8D149+OAPx+SHxC//JsA360m
FxeP3tpaKXAimb/9PkBvrbRxGj+iTWarBr+C4wrSOibj81zcwAW1e23B2UpiHV3QCkO+4g2Eo9zl
/UBCTjAQTmMYDj/nvVikgCBJ/l4lZwrdCLQicDSSGmz857csc1he4nepJirVtKcUzf//JXiZmHQI
qfSNzTM2ZsDdQldCkndtlpE+YLR4zRw3Y1wpi5n9lntdjWnztNBic+8d0+bgk1U2M9khjuxS1EIg
SLyJCWGspisISZ+e5TS8eU3Uuf9lj0UKVsNGHky96K14sTR81n3/yp5MwCy3s2bIw0/fdyvQ2pEQ
gE4c126C16Fno976g+H5UPkplbrKMRO3JY7N/8+dYcXPDNWZ53kSGUDOkAreV2CjEce/YWmeTIji
PDOvc944AcaTlk/UDkgYAUVJihK2I9c=
`pragma protect end_protected
